PK   �x�V*�ŀ�+  �3    cirkitFile.json�}]�丑�_i��K�@R$E�����x��>L7�t约�oV֌g��/�̬�Ee(㨫o��Jd�(F���ծ��y\W�]����=m�����ܭ>�������n�y��o���?���������$�)�r��u��en�Dk��L��&�I�*-]�ʶI�b-V��xw�ɖ ֒��+A�W�X�l\	b����ڰ1p%��ec�J댍�+A�W�X�l\	�G�%[�Gp�|_)�Β-£�K����0�"<
��d��(�N�-£�M����8�"<
��d���w�Ex|���Q M��T|���Q�}'[�G���l�w�Ex|���Q�}'[�G�������_�]�+6��|�y�P�6�_}�'/�UX������yܯMդ�U6iKQ%:u.)��I^�,�����`H��s�XI�I���M���.e����2�)3)�����$��l9�	L���xz���Xt��cu������Xtb�bu�buE'���Zcu������Xtbm��3X�A�I,:��X�Y��tccj�S%Ea���}�QU��պDJ��v�j]ƌx$���:ê=ê�Nbщ����auE'���:��.���Nb�u���:���0���,��C'&����Hpn"��	������'(X|��[����`�I0�na�?p���'���%E����
���C��gX|��[���y`�I0�n���7����&1��}6_gI^
�Y�L�T�Y�V�rp�~NdV��(�b�)y��ir�Ә�
��qUՅț"��O�΍K��u"k�l�Z�䆽.��	S�i8y�	ɘ�2�N*��Z��J[��Z��2�e���̘���P �G��s-�2c�O���ڴM�*����&E��I�6M�����[=8M?'�� S}a�J���<��Y孾vI�dݦFۺ,�V���O�Ƀ��� ���)y���4���ɡ
���[��2�4���y�
�#���zpJ~SU��T)������l�iLUMd�7�H�a6#['��@�������[�
��f��x�Y}�U}f���Շ��g�U�5��[�L$Ýݳ���>�iN�m�3��SϬ>�=ט��Ar��$G��I����z5����gv��0���L�`ͭϴ�������1 f���,�Nͭ�#�I��`A7�=�R��mY�6�w3{[d��ԃ�d9�G�������x'�y��4��U�9Q7�H['&K}�k�'�L��5M杋���T�|s�ys�؈��y���Ķ$$1GU#�º$�3�+7m�7�H*S)g�����i?�Hofi?�H���z< ��6noev׀�an���N�Ulx���w[ֻ�0��0��r��`�9�^��<7Kʼ��LaH���sL8���ԥ�򤴭��.DRVZ'ua�,-
'�v"� U�;.?,��9�TBz%6�I����ƚR���Ӊ���3�����q�I�O�I��9|jʦ�|H^�ʧR����IU۔���%��KR���I��'U�k���p���t7���<��8���xb�Vu�
��E�G#��-�&K�K��P�m���z�I�����ͬ�E����.)u]'Ejt]ɬh����q��L��D��a��qF���H��)1�d�Pi���lƛcт-m^;c|��z�k�")�.n�*��(�	['U��:�z��I��N�|���C��/��֔Q��w�	�PF�\&I�
q��c9�լ�AƼqG�2�-�v�3���J�$�Ab�wģ<-�NDBt�Naf��0(�
m� �K,Ŵ\����v��ַ�lWT"1�%�6eYL�ˤ�qE��Ǉ_R���K�5I��&�z<�$U�������mR�~v���~GO_m�;>=�������]�D	���1�@�z�z"�����$���� 	�I�1�@�z�{"��� �$���� 	���1�@�T� ���8����Q��� L0�-a�%�@������Q�d� L0.aN%�@����
��Q�$� L��������q���?̏+�GI:\ ���
��Q���0������$�a(/��o�R�cs������!M?kH��i�!
BjH��
���å��֐���!�	\*P�K`��1�����֐���!�\*P�K`y�1R����bE�K`���R�z]kH�����.��%��`40$�K�u	��e�>Lb�b���hG. )a��k��k��k��+��ǋE�v��k�#���"u�L��ڑ;
�b��]&[���x�H�.��-�v�n�X�n�@;r�H	�$c�� %,��-�v�N�X�n�I�A;r_f�&�[ ��eҲEЎ\��\	[��U %���n��@JX&/[�ȕ �.�"�В�2yY@���2y�Z�X�n�L��e��h�H�.�����l��l-@	��e?H���e�hJX&/8�A�]&/EP�2yY@���2y�(Z�����y�n�@;B�?�v�A������!R"���2�B���F�)%�'y�i�ȾߙR";ugJ�쭝ku ��R��[���|mᔭ8b0�;j5WƂc����p���\1+�Ι+�V��:-9b0V|:h�ڜӧgC�6�E��[qn]�8���Mdui8b�V\4Y�u1V�^�b*�:@
KߡL[�:�_*_zg�B�5C�ը��[��C��Ls�:�k[�R��%*�8@���L2���������b�5GN��v�dZ�鏢��Ow*��t���vO�T��i7Ce˞�D����mD忞�B��H�`�گ��� )Ws*S��*a6@��6��g�\m#*��t�I�Ş�TJ�i/Ee����� �jKS)�R�~�� ��R�R��*�5@�հ�Jm=�TPi��*���Q��R��.��zZ
��zz��,=�w����~���<��J�<=mAeU����$_��� ��d6�ax����� )�c)"��v�̼�X�� )W��� ��K%�H�:�R�|R�N,Q�}_����>�}��}l������m�� A~_"���/HЁ��$���At��� 	:��B��}!�@���D A~_"��#�/�E�6�m����9n��#�/�wK��FI:��b0����9p��#�/̇K�GI:��b0�����q��#�/.���0?�`~%������
��Q����L0?�`~%������
��c� ��h���� �#��h�0�#��h�@�.�u������0Z*P�K`���h 8��
��XG�}!�����~_��C�h�@�.�u�����@0Z*P�K`���h 8��
��XG�}!�����~_��C�h�@�.�u���/�p����~��k�c��p�H�.�v-�w���p�H�.�z-�v��.��eүEЎ����"u�L
��1~_�X�n�I�A;�����2��"h��}�b��]&[��/\,R�ˤd������E�v��l�c��p�ȕ�e�EЎ����"u�L^��1~_�X�nZ[&/s�b��]&/[��/\,R���e������E�v��l�c��p�H�.��-�v��.��e�EЎ����"u�L^��1~_�X�n���Hho���K��征ߗ/%�_�~_��Ȟ��}�R"�~o���K�쭽�� c��C`����`8v:�~_��ǎ����z+������ cű�&����`�8v�~_���+N�Z1�ߗ/��j�"���\�Nd~_�������˗r�+��}V2^��^�j��� 1����}'Ő�}�R�67�ߗ/����}�R�~�ߗ/��v���|)W{5��wR
�ߗ/�j��}�R���ߗ/�^����R���|)W����;���|)W����˗r�v���|)W��ߗ/�j�K���K�j/d~_����K����B���K��2���8M���K�Q�}�R�GAT~_��^���ӑ�ߗ/�z,E����B���K��Ed~_����K���K�:�}�R���d~_��������ܯ���v����\�W�n��f�<�??US�7���nv��?��X��$Q�ns�J�8o���X.^��6�I�8Z�����!�A�aH���5/GDK�ֆn��i ���M:�0��h/m���o�!aS8EZ��],$)	�J�c&����Mp^-y{-8�f޿�yu��G�~�ȫ����-Λ#7���8�rzZ@��f!P@>���@�^�p/�ψ�C,5ɯ�d�8{	�%�z�д�EhJ+����e?�T���%kB 2�'�9���srv�KB����Z M��zp$��!N�3dx֟3��l�ͣ����=h�<())"�ұ69s^-�Z�8-pmÐl��(�ٱ�ys���|9�sz�����p�	��[��\6q;#�EDM��m��n�{w$���������xZ��5?mn�u�X�-���1��
����, ̅>> �z��7^������^\�� �M=ķ[��y4���&��C}um8���m9���Š��Z�z�ڿ���4�5B8��\(_�<n�_b�<��b6���|@��|> �>wq������G�]�D�%�f> n���Ul��f?�AFRs�� �H? �b�"�DO6��M�3z��6I�}; ��# ���kދ8ܾb 8�?f�W�EI()>�=w_ͼi�-�~m3�#[��8���� �-�\K��b��$�7ٿo���3��I�]��7�����=jGl��������?���m�|;����rS�����P��0��BZ	�Stz��-6�����N"�"�G�лH��ЛI'}�=�| ̭��yy��I@o�є�ߔ���o4�ݧ �M�����!X��y�]?�}�z����m�����yS������r�u��e�U^���\�/B�,MLl�gyb�`�=K[��Y��(�"D�R�D�!z�+&
�ѳd1Q�E��e���-B�,]Ll�@�u[�p� �)�/C�8 >T�(_�8p�sq ��8R�q�ۈ��K%���e���J\ � ��/C�w��@ģ���O���e��U\ � ��/C.��� �S�|�pM��*�?e�7��_��̉���^ 7a8�^17D^A��s�r��ٖr�%/�1���'�
�?�_����)X)XX|��k��j��4XX|�O�X�?,>	�'��wHy���'sqW�3�:3�:��$�X;��XX|�O�s��r����$_7Վ����� cJ4�n� �CxR�J�i�D�%���J4�ny�CtrF(���%��	
�D#���:D')`���[�C����J4�n9�CtvF(���T��
�D#3sz�=��NZB�@��Ylt�2<H�s�X� �j ��9A'5!`�@�J��a��ǤP����:�\
���
q)�Rt�F�{
T���cT�΀�/na�� ���cj ����@'D�C��J�����`�����$0�1){���`���Ґ�!P)�J��S���+ٓ��r��|09H�3���`��\2f�`��������lUӛ�fS����+�g����&���bΧ�c
����TaE�_h���r�+�k�Ṓ��V������b\;=�?�$bi��
=��/���>�y`>���ǵ�~����dyy(/�VLi�6�N�8�` �`�Y?�b1�g"�I`���(L���@Gd��E��$n����O����ٶ�5���\#�r��ѩ�)T�N�7�Q�6O�7��H"+��ɝٜB��f3QÙ\��4Y����^\!���:��fiQ8Q�SC��Do#^����}�Dg'^U��?��/��'2���O��wϫ?�"�(5�$2�N�t�f����<c�K��V�N���io,���R��8a���N�?�ؤ���zVע�.�[�6�KJ]�I�]W2+Z�&���~R}.�	c%՟p��΂Tb�'՟N���Ā�IM[li���Ðֻ"[IQw��ު�[-�r�:I�'��T�:I�'��H�J�� r�N/��&$�^9�M�<�Kh6A4uJ�HZM��%ҜO�g�f~��c6�y�:�M�M�ޥ8��xz��LqS���yz��U��3SV>��ze�&qE%��ZnkS��d�N�?�9��>�T���O�Ȥ�#2��ĈL�?1"��OL����~�[��������R&PW�\uηs"]��kg�]?�F�n���_�Q{/ݻ��I�]��}���~���>�C�~ư���>���d���~���sP]������ǻe>
߿�2g��N_�2�p	�W��\�����U�P��P@U���|��J��K��h�<��1&�vZ�ݛ}IJRh�����#����{;!ҽhJ,8�FJ�|'%�}e��F�JGE��3{>���f߹������D޾���gH���p�{�p�[t�V7e�]��� ��4�����3tor[S��r�ysS�.�tj�-N�Aý�)@�s�{���\;B����or�S�N��yT������A�b��Mn�
��|�����t_�ƨ M̷���Q������t1��%n��Q���K�0��y���m* s�oq�T .��B����/r#U�&����T��_�27Upb��K�Z����/q���ʾ��~�P��C7�"�V�Wi��>x"��d�H��Qz|�������#>��G6|�e�#w|��G��Q<�'m�P�E�>�I2T�<)D��'��P%��D�t"C�ȓRd�yҊ�"Oj��^�I/*ԋ:�E�zQ/v�E���B���^T�uҋ
��NzQ�^�I/*ԋ:�����M��>���<�����i����S�U"3Yw!�KJ՚����v���ڦk��?����_�~h�}7�I�Rq��(qo�A�tm��7y�2D"�E/����ž���������f��4���O���뼕W��~�y������߻�w�������^c�6z~�x�+��ӧ�/�=���]�o����?|jv�<mʇ��o���=ovM�z���}c�T<>�E��5�) ��ΐ�� �P|���o�^?&�r����dvo�
;T���+�֥�~2�ǓL���ǥe����L뮯l���cu�CZӻ[mw�F������S��Uͱ�<(���9+>��_Ru��<"ΞXw��f�O��}�D��b�bƝ?��O�������@՝�S���ȃ,V��jh_��e�~�gO|�>�ŝ?��Oze�~Q��/���A3�_��{�Ĝ?IOO>��������s�����=Z^���x?����>"ɭ�
�����?�y~�wT�Aj'r��ݥ��EzG~�w�unU�m��e���eu�M�(kE�D��~��E�%�S���zR{fJ�������Y���7���W`/�V��y���c���i�ওis��pJ�,'�=��e�q��vj]+��iR��_��Ju��4�i��⠻�!m �N����A8o,Y�^<j+ƞ�b0���pb�Ҿ����*�^�<U�H��,�kʤr&�2�,)�,|���EZg�Ɔj"m��i����}��t?0J)�n����j��mj�G�C���W5�X0�O3�F����
j�����;LR?�tR����N���@?� ���W]qwԕ�vS�������D�:�"�w����*ߕͻ�_�ϟ���~��x��?5�w}Xz�����������|'|�������E����޴m��/x��_:C8MҜ�}��޳�w[	&����V����N����?7�O߿����єE����Ϗ����s�
fX�U�h���Z���Eu��c/9�zy���Mı�>=C}�Ө������7�R_�bW�E%�A����w�ݻ�4�L�x&)���٦�~x����w�I�5�qҏ��]��iV�*)�<OjYj�j\�۶(t�Y%���S6S]w�������0��c��������ܽ6R	i�)�����:����Y���k9��T߶u��k���M�Ԥ���(O��^���ٝO�/&,d���^�Fe���p|�r��*?��{�T��ß���aŏ�ʹ��n��O����vZ�϶D�_*���]��Ff�_X���R�;�u�G��kO߬﴾7}��^�r�t�2q���X�7ܱ���0]�#3���s�vF�x{�;��˼���c}�����.w���U-���=5�/�hN��M0^� M����h1�c�'�dʌ�ư?���^w�l>��Q�MT�1_-��l����w���y��6OK��6��a�#�#��|�0��\������'�L�n��
�Adf�Κ}r��!&wy*Q'ҵݺe�U�V�զ���[Q�/io�P����@Ə~�������5��2�{��e�r���<�k������T�ަҨ4?+e}|����+C�;cSeNN�{.����>_��_u������_<�/��{!����5�iՇ�:�@�����9;.Ħ��we�w�B�w�,�3+�q�7�>�}Ի��+��47N���M２�s>]:��;�M-۲ەSv�&>8˒ԷrⲶl���i^΀���2��n��|��c��i����|�G��ѲS�p6�fm\&N6����Ѽ�,O��U}>�H�F�$M}�ZI�ڧŉ�!�m��.K=Ti��P}ǅ��񩽏��px�x>4��{��g�P���X/�kU���|t�����k\�>�I����'۪�4�ڤ�9U��ZzW�r���++W�K���|}��Pˤ$G-u?��C�N!�}����7y��6O��3R�"G G'rV�l��n?w����(y���g��k�WS�7q��{�a���O'��ntu�����>��O�Rッ�-�Ĥ�׼)�i���L'QS��Y��[�����k�P]@g\�����|�+�)�u����ݺ��[�����J����lG������i���Ku6Ԉ��Ag-kW�|R��c5�~.��d��a���)�y1���Bر��ͳ�I|B�ż����S�Z��Dn*���N����V#��A�C2�'�D/�ҹ*����G+?E��k��gn�^�f\��a�)�L�u���h��|:V�q�co������h��G�-�o~���$��5���VY}��d-�>��D����(�=Fi!�Z&M�;K-+����_UV��H�&��H�%	A�T���,�i?���~��i���~f���/���DW�i�OR�p2�pA�ҊST��Ɇ�Nߜ2�uf��9@��S!Kj�*)}�eSmeDUj�`������y�;)��Y��V#�:g;���e1�� #�t�;̌I}���އ�~,?�1}��3��x˳�׶ME��§O��uc��)��4)�Bu��Uo���y?����O���>�Pvqז�[%�ک}���g��0|ZrP�]?]-��W�u������']�y�UUN6m�V�(�vB�' ى�w":]?*�ދ\z�0����t{���@�[��U(w��}�׃����|8���_6��S7������;c���ӳ�6)�����?�ʿ^����(�OM�Ǘ-�����׿m�_�ӷZ��������v�a��C���U���������<~[��n>d�k�Q�3��]��H�^޿/���v�����e���ÇU�C������}�}�������	_�����g�n]���b�0�Ŕ��X��J�d���X����ƾ���1���yg�1�����ζ1G���b�"Y��ˆ�x������D\3'x�}��i`J_i��"��ӑJ�q6xcXjܸ��yc1�"���׍#�иƝװ�7��/�-�\cX�f�˦�*��qV��8w���g�">���q"t��kuj1��Rl�X���2Fy���qV�1���k�gSj]K�Ϊ��s����2�7�E�3� �B��<�n(�H�@�7���1o��i�#pg{ƋI��g��<M�z��ss:3ځ͒�Q���� sX�&�q.S8i=b�Z�M��f��*�kK��� (����:�n(���7q�n)��qs��S�B���
�R���M^	o�7��%��q۸T�M�.��.���Ƌ��V�d�m�8;�h��C�H�fG6#��A19�?����c�n)�G�#��
�bAG �4VBl�'o�f`E�#p����3���4K���/7�I�f�sRc
�%�o])��i���2w93�mkoGZ)���2ym�l�v*媼�FsS��\Rt4w%u�	s�Fsv�Z�iuK1)}F�����vP���lf��#8)$�PO%�-�݄�����T/;�ͤ���"n0L+��!��޶r;kĤqcGL{�9+r��;{��es��t�7ȟs�r�PJ�aj��Cc����3��"��4�h�=�7��X��8w�=���G��m��x�.�-���ѵ9t�OM틚�5������&x�7>iҔ�Xd�D�TL�X9y[9E��2�����O���f`E����wݵ��-3�������"�-��i��X{47Ƈ3�"�q�l{,���q8�G-g"��-Ũq�i�ZS�@h�7��Y�et���0��@7w����X��Aȋ��=[/��	u9�K,&�w��qE�9�^؟�W���ר�9��̽�l�W���1-2֜Z�Tl|��㾩�����C��ؒuFJf�#Z�ؐv�p,^�B��P���G�ε�j�H3ލ��؄#�e��>�D^f����s���׭�g3��q��2�Lm���[�Q����:�;����Y^g�e���a�0��� �Xԥ�7���:-��g�-r�����g�-r3��?7(/�yl�lP�ر}A�ع�P�����6Pb�4�|��R,�g�H�6ip���h�4����o�U��Ŭ�X�G���_J�Ե��Ό��N$��\�vv:\ϭ+���c����C�ٕ����c�Q;�,�#�斉��9�1���|^o��h7����k4�y�[�kxƔp�o|��f�y���-/���2�VSt7wQz��8���f@CY�M>錰&n5�e�h�58�L*4�[{��<��P˜���E�K��쯣��<<|��G�ov���i��3ɧ���7������?}�o~z��������PK   �x�Vs�7+5J  dK  /   images/6c71542d-16cb-4630-930f-71c4de5e1144.png4�4\�����G%�F���w� zｷ�e�D	QB�����+��=z������]ks������s�Q�*�xؔ� O^NJ��|��` �_Q3?� y)q���m>�Գ�LWm�5��G8�� ��0P�����h(_׎��hx���๓}��2�Y2���e�`e�e���Kw*�/��|b��G��,�\*k���-/X�F��fg��œr�z�cvvJFK�G/�/i�)m�b]��8�X
�LTjYx�*?>��98����O"2����.d+E]r���q��JW���5,�3E�G\w���_����� �Bĺ9���� !A���7�D�L�2`qx�^2b��z�-|�_�Q��o���O���|�w��o2r|u��؁�P,$,��~��v�7�5==�ʕ�����I���1�B'x��G��'�w��*��#N����G�vW�)�S�J�К�V�%�0�=^뽌�S�13�E�j�^Tj�i�xJ,_3��������T��ٞ�Rd#%*1]{<�+KSH�������`)\�}�^�X&.�.C�f"��#Dj@���a!�B��L ����ecŇ�X�\_@買Ox��-�C�����?����dʲ�J�qQ��s�JC�е9���tx,xXb60u	Ȳ�l�Lˢ�:�l
�Ð��ق��}ǿ��Yn�x�t�E^�M��x��-G���M��άG8�jε�:��C��#�,t�H�M�Q~O���Q�)��%#�!���2�cS�!)�����k�l&m��%�� X�)�t�琰X2�_�N��DE��W�������(�]����R��TI��F���Q��A	�
��)�)/L�<�٣�п��yR6��n)R���D'�-�G\
���FF�K�Ă@g0�/"��9�	�M�#'�9H�a�
B�X
w>KF�"	�|s��/iIġA���a>)5�:뿦���[:y"�B"����N���/$5vq!��}�Y$>��X�3�CF1�y��h9�T#���!� h��+����ގ\WggЙ^�E�-����]�ȂrO�Q�����#���:NSA�Q���|Y�,	�����Rj��[�W����vHpc�z/�4g<QZ�v����&�^�Vɭ���a#���(�|�D�<��MQ�KO�Ѝp�/ �l����Ѝ �d+��ྉG�O��Q��{��ڣ��u6\�@B@����0�g���㒒��QF��c��
MHBQO��3�V3�rP�� ����V��J$���fvf�����v�Y{�{~�Ű?�������E>�=d
�=hh����I���Ě��$�/����š�6�:k��D�0�U;��`�e��gV71"�qq���O�,�ظ������;َۖ�E#�3�=乚����ԭ9LZ?�˾nP�6��e=F@$���'�����`B1@���a��C��4	M(���g�1�Kq��t�-_��,����pV��7$��铂��u��)��eɌ����=���m�������II(8=33�Q~�˼F�~�/�g�K�PxPI��y�6n5[���i���X�O����ߑ'���'�à� �����3V �
��F$j�ö}&=�e(!��s��M���&8���(Rjal#Pi�4���O�>%�|�jm��7o�s۶|�-��w�}�7���aގ9��xh�r-�H�L����=<ʪ
@BD�j�C�r޾�5ȱNw�#[�S>Y�b�I��������V��[���|�b�����=_�kX�Á��FpI�����V-��-y��B����D����^L�4-�G*L����pz�1��
U{�^��6)#g_L��B��['�D�Li:�aAU��ɚ�I�I+@����ދ�4��ޑ�-��؎��M��L|A��"�É������ҧ��T���}*�#O֪�x���ٿZYZ�>�$�������~�<lc�w���]��TW�Z^N0�ZZ2�̇ȧ*�p����;Sc***:����hkk��^��?�%T[��;Ș�������k��g2*Q�����I�ʲ�I�H�(�D��mN����7���X�j����M������(���Qn4t��Q�����}���������@�?�̉������;��&�wڷ�����ɰ�I�m$���2*ʠ�:�Zh=�MX���e&���C��X7 �Kz�G���O#����６|���������m/?��l�"�
tIr���$=�е����_��m���C��^Ӷz6��+^���-G ���%�"O���_鱧%��ώ9��r�!����d�; I���|8˗�(���8���EF��׎W{>��Ńl2#֏{��^szdM�FD'1i��	j�V>�*)Y��yq1��8�	��?I�Qz�C$:��h?�􉅲�_vb/�� b?��m	8*�䍳-������@�{��z���ͪdԹ].��;{���X/V��_�*b8OP�(j������̱K�w܌t�Hjz�:�����Ҧ�5�m9���O��Z=,��X��\�����}�W)m�����CKPe�PS"�N��Jq?WgG�v��kt^E�} ̩����$�R�t_2��QRRv���!tZ[G'x�G���| � ����˥֝�ʳ/5���XP��R�/x(&�ݟ� ��xJͣٴ�[?n�|��ܪ������l�bZ���;o(�5tx�b�x3k��I�Q��U��c	GD'���!F"�Є ������}���8��BP����4f9e[w�o��@�l�&��E�1��p�˷�HQA�ֲP��S��P���n�"%R�Q��\ڐ	(��ۘy��3������Ue;�?�u��)�-p1w�s�Dh~�	���:��;J�VF,FR�}�B�.��Z�Q�g�9���O��!Mr5^Х*V�غq�}�g������d~�xA]����H��ː��w�Nf2 c����R��l����m��]���oyےV�:���i5��D9�1@IYy���X{��>ӹ*����D|��w��¾6}k]�5a߾PI>!�(��B�d�jg��/��P�U��\���l�!v-���1�~�{	C�����7�tp��ফ���T�|P��?�DL���QSS��8bBt嶫������~�������*��[�8]�Ă���$���[m'��4�:i��zP�$E�o�/�2&�������Х�'��:E��,�������l��H���g����=�*������3ܹ`J�`�5'���cD�rN�k`��[L�p��& �S�kV�g��� ]��^Xˠ�;�#��G����4;<��ߗ. ���\ 4W�	����2K�n��vd�L.��x�����e1lC�~	vjЦe'A>s�����%��X������	�+�`������S�8q�Ý~�tgc�܎묎�������[��?����OMu`���3�tߑ��v��۷M����}*�3��Z����K��n��9��d1��>6a����\���YZb�Y�閙�%�2��td*���%��p鈈Q/�����R�_j�HQ��%����k�`�Xo'�VͶ�Gn�;:�+kD�<=�̬�`Lj*���&➞~���lUW� ����4��������*�2����m�������vH��"
��UI!e�N�<"ȇوHq�^��UduW+}/	yo�C.A ��ل(AS�
���+���h���J���}�vCF�!ԓ�H�a�ޤ�;����HRS�уC7���rMC��a@F�,��@urzH��Z/�Ns�gK\ۇ˵�.v����/�4 n�pr&&��DP<�<�
�e���5FO���3UТW��U�~�m��� m`*������z�eˣ�g�>�GF�1	w����o���smJ�M��"�?o�u&T��2&�OؘT~_�=�>s�Lo��K)�<��{ӱk�baB ��TC{���o�B@}�ıi���@�FEa��Q V��ؓ��f`�G'&�LMQ�HOO���`���.�é����F͹�F���F)ju_6��4,P�<!A�e�2���m�Ȼq����4e�����%	MM �� �&�Qr�G:�ذژD�K��@G�ϝ�R�u�+@�#�i��b���Kf�f��M��[����=���q.Ȭ��z�y���9tU�d\ò��pi�xAj��-@�'ڟ'f�	������g#m>���J(�P�:��� '�p�bJ��$�9��v���I�(�����ųv�w�^w�77��1�(��Ǉ�������ՋY#r�J^� �����B*cTlB���
����7n����_�?�;oOM�
|8�ո�������BWM'2�bآ�l�C���+Ε���|�����H ؎������X;ݷx�.L���S.@-V{"L��!���+�ao愯i̹(ҋ����F���!T��z���<�l\U��?�� &	����7s�	�'[[[+�(�N���Kآ(9ݣ5n�|�����ݍ�F�o4nXё�̩�JJ�6�pL�I)����-﹠o���ѿ�ҋР�]w���]�oxx���΅b��w�Q��\`��5^�lu;�m�]��nr�������|g#u5���J�|��*7�\^�4	������ Ȳ��_�)��lO$�=�>��3�q$����������9��ZT�Z������^h�?�pV ��uϝc9f�铀IA�#�� �<J"_��"V�L{Է�o��6"t�A'z�#�}}j�Y4�&���,����Ö�Z�rLB�t�;��r�m��� ��4d�����>i ^d�{�}���H��!]E�Y���]�499���x���g�2�����H� t
y�f ������:��Z��3%"
�L�����>i�>�T����������5������I�����������T�Rl�i� �N���W�0 :�jjL [z�&! �Wt<�ӊ��M8�"m$����g}�@�d��N�?�:�	�2��p�~3�=K!�S4?����giee����wfQ޼u�Vi���l�3�Q^'�X�r��PN���F�ÁE՜�z��@h����v\ta�:��RaȐ�V��Ac���*�'��q�l�d���l����2�*�����}���J����(���dA�镑L�F��-u��	OX����,���ud%#�x
��s+b-'�tr7S)�O%V@i��,�3a�;�ĺ�S�����rCRGa�klW���$�5~|wY��o���}}��y8wI���P��e���;��o�,�7K�Z:n��D�UZ�Q�ܾ�|*7��1k ���@z�6 �'I���a�3��ˁ�p�0���56���|��	�G��f|�Ώ�3�;���s��}1*�sZ�䦘����rJ����F%��960|Ռ!�.��� \J�wv	��Gq�=B��ڕ��$i%+��#�����N�dR$
���JJ$��g]�?z����)o�����u�ou(&�u�����t��^(M�:���gֶ#��
dW��Cǃ�b��z&�������l���&i�����dɎ2��MQ��//XT�p�7�2�Ka�Q��4_���hblPmCCC����9e���t7��G ������A���;OЋW���X#ڎi�ǧ�J,��_?�V�<�D|�'�����v�x������/��� ��9����B�Gd��O�C��^���İÓ�k./��M<�8��w��yPp��`.��A;]�������dnY�fk�Z���-�tŭ�߻zX���j0;5;;�ے���vʺ�^��Zߘ�Y�e��b�b[���6���;�u�j||���3pq2h���<7%�Z,����籝����~��R�p��(txyŔ��C�j$j(����Q�t���Na�?�|NM���5_��U*:X��@�c�#7����{	�H5��T��������:i�M�����%{<ʒ\RU�a{�0jj)�,�*�^`�^�b�S�	������W�>�P������n���o�?�;5����G��l_�m�[���2��iii9Jf��])�ÈH{�S|ŵL"^�vtKZ����ﾱ�,?z#��揞�V xŗT�Sm1��r�+E���B��I�E�/�[�����.%���QLw����V��g�{�-�>�k ����=���;��^�cit3Ӽv=:j7�[���q��MVK��Q�I����*ݶU�w ��H�G��4�^K�Y �0�]��8J�z�kɪ)��6j�N�Rl�6�5��y曫Uf׿v�L���x6:4��Q��~������P}����Co��<�6~Jg���ĒF���/�?v����|U(K�����2"bʑ׻���cJ<�0!���fl|�+�I?��\rc��?*Fb��q�i8�iY:������q4ug��c �ɛ��g��PSQ���ճ�j������.1*.:J3���H��.�����%S�[�O��p��i�f�U���l\�������� ��p/p��6tHי�+��!F��9hu����x@G�T��ళw�5�� P(]��0�����6_x��XʞN�\V�:aX��|il��3�<}�ҨOyO�ak(K�`6:l�GZR�G3��(`���'q~�/ϰ,X�����n��Z�m��-�F�Cf'��i	��Q���g�����Z��PYM:������o�
a!���Xt%Ҍ�Y�R|
� � \�����D�_� �8�j�N��jt�迟M(!��S���cn�x��T��Y�V[3�[bƗ��R���^&~~����.���n�.��&���Y��ZM�e�q[�&gb�p_�z���{:��l�K�I�g�x_K�?w���4CÈ9LW�غx]��B-t��ז4�)��g��  T�II�@1sX�?�To���Կ�2���cOլ��$��U�&��e=v�5�K>;7H���~*�j��p᪴,n�o� ���w}:��YD(����J��Ƌu��l�*=�lښ�1q��&"��@B�͋�J�2{A KC w���U9�,9�X�$�����,���!���Ð�ȵ;�]��`O#�$�	\��oJ�	Uy����N��G��.�f�P6�GFy%4=>��_ez������E�m��K�KV�d�MnV������E���Ӎ��
��3�]w�:�g��d�Fv���7�d�+A��OfC�DD�z����ĸ� �`�xj�B��v�����H �O�BAv�zd1J�[�Ĉ�0�]�l�~���3F�0�H1��Ԯ���W{v��d�T�
�V�$#�M,,��d��(����lwƐ�*���Z#��������y�4�rؗg�ۣ~u:�۳�y�m]��2�`�z_��Ȃ��r�ni�����7J�Z�t���}����q���#~�z�:V�ʦ+�����3����
j@�c�t�r�o߾537��� R��'Q�Q��?��dLT
�opJV)rY��t����=�K�;ep4_¢C	rz�\���}e����1=u����V�����x͍�<�0j�:HH�D^�BaHj*�����A�r���7:���߶�$7�g��������=�=Ze�:Sy�j���h�s�(9hΣL�gJ��ͣ�K@��K�i���+���IBUm-0� I�<�Uʟ/�~Y�f���c0+�m}�ݵ��h���r��� �bQ���P�`h����&�72�_�6V�~��J�Z.#L������b!	Ck��?��7���T�Cub��ag���<>����Β�_�ڋ�|j;Q%��Q��lN/q��4S�^��������^ ���Z�^�|�H���䐇����	��@���8�����O�@��\1��_�֏7�q�p{�PH7�'����͍�Y�n�l��LF�����+���3�G6���c���#/�(0[���t���nZՊ.�՞@�Ej�Ɔ9	�5=@� p][+[cY>��B3�]����$!Ќ�h10m�1�T�c�OY�@A}�-1������^{+���|�j	���N��w����Qm��{�M��<��c�w�G�����������yCG��J+1%Xv�L�N�6p�����H�����>j��l��I�2P�_l!�G�zz�9u\��������)�r��`K@֪�+T_�$������#H=H��%C666�����*�ХeP�D	�xW��V�f��� }���ng�Y�Dic�8����� $M�x� ������ɂ�{�?�{�M����t�&'U�c:����JS�q�^�O�,x�#��
���h�������C���%�WX�6���{���s�Y�Θ쌊��:i.�ä������NJ$�HtX����q�*��>�NI�����6VH&1d���PRr�CrT�&��U�?5e��D�~#�|lm_�i݊�Z��x�A4�RU6�L��PLe�=M2Е�6]߀:W%e_5���ȼH�L����V�`+�:h�@�ϙ�vZ8�kk�Gal#��D�������.�?�?���� ��gӟ�����
�t�9��_�%1������9kʐ��ߞ��Bm��B����0P@H2�|�,��i��[�?o/�H���P����:��Th_�E*��H��:Gw��������l�
�fl/�c�����W>��~]�v�ӳ��>ߌ�
{���[q�~l�I�՛p�Շ�k�Bov�JP���4� Bh�;MO����������c�($����{D��������oo>���:�����#�1a��r�����M��G���8��`΁�U~|́�lp��)�q?C�cbf�jm-�r�IR5�����u�ad�1%xU���;���>< ���װ�)x�viG�5�P��ȗ��c�S�q����\�t_�_\���9v�9���$��	�7:��?�,�
ݖɍ;��UJF�Nu�](��-��'7{f�ֈ*�uI���yŤ`�c�/]@d�ԭ��[�h(
�ޖ`��`;�Mz�������xL�>z�ߎЭ0Hh>4��~7�qZ
	F������dx����Bm�ea�j��f�#��)�sU�?諔$u�H���py�b��
�ߧ� H���4R�a7�13$�(s���φ<g�;���Ҝi��@��F�·�'G2�K�Ee�aL�Vԫ��q�� 4���e$��ϴz�s?ap��!�&�ρ{�o%*ɗ�ڭ��qli�? 4�}�*�������[#in�9�D��)���n��li�{{0Zځ��s�֋_z��&�	ӟ�Hݲ�*��F��U���0}'�%%W[�y|��gKf�9G�Ht6P��`��{g�z���&75�8�.�H%e5hn�r�f���f�3i(���E�T�BW��#l����?4^�5��l���B��p��n1H<<����p 4���v�"w#0���4�7{>�1{�j���cs'��I�~��*�F�,m�А�Cԙ��u�Xp�C��
���jʓ����T��6xs�X� g�� О�4����X;oP����u~s���`ݲ����^�Y�c��@�y!���GP^�\rXF��B�+C0Ȝ[�)j�|�q/�ە'�%A o���I�g��Y��VU˴�`�%��%.��0ժl2h��P�R����ro�Qo&n�_+�}������U��G~�,����kzv��ȡL�?Ǡ���7�T�v�N�/�����&��j��p�Y�k/�7{�;�R�T�Y�rA��r�pp�Io:Ͼ2:�w���hm���A�BZͻ��a�Y���^_Ћ<-i��]���s{(س`Jn��P�B��~d�[i�Z��P���˞ж���q1���g�c��*gXQ��X�gϤ�2b� ���8�<B^Zp�iQ���4	N�|�5b�2Ijel�W��P҄����3a�hfP�NL�;��{�n"��f�ΤB-PE��V�ދ
��y�X-Y�l���ڎz�]N�7<���v�n�ta�ڃ�5���M+����&\i^,S� ч��`��C�Op����V�b|��7nXuL_���d���;���������_
�}`#������<OH��0�$�u|��$�Ўc��� <`��h��,�is�5��q�#����?��Gm䊊��F���W:Q�^�:[�`B�J�Vw�f�I�ƛJ̋�<W�ͤ�6e�{����{cƸQ��2��|�G��]����h��síp�DsD���ؾ�nw�՞����NZbؖHZ�v�W7&ڙ;wB˴-Tv�8�m�u���-VL&o�g=�":��+Z�
Y��$Q���cF���`=,�$��:_���(;C��%�6Y��B��%-�k�=z�}���~�%̹F�/6� �Z�d�ɬ\��?)O�����A&>u翃�����~D��>��Aƺu~�����ľ�6��e~���v�qJ�r�L�
҂Q؍�G3��`���ц���iK�|K�����w�����_�-��r�v=4��~Ŕg�1C�\j*�|=ެ���~�aB@�q�:�w�!�p��u�����Z1I�0��|q8T*�y!T�>n"��l���Uѷo.�c=F(�s�-�L�[�x����)L5e*��l"A��j���t�QE��ԑ��,�LQ�Ӆ����풆��w�6pn�_���!#"�.y��i�i���Fe/��,L��)�����Zef�a��M��?��$��.�?�p(p8�ej�=�V�t+��+�f�+ �����"�u�`�yM~�/[{��٢�]�^#��6�{�w����c��0JJ	�������qn��.���@}p�L�AV��O�g��4*�Ǿ*�� )9�G[?S���
c��ޯ1�ӨW&{��Z)�D(gH(1r|�(�^�<�����v*��4��j��i�F���\(����t�5��վj���$#�ԋs���@��&��������ٳ$�`N�%�`.Q
�d�VT������/�*�:��-�vۙ��K�f�X�/Gт���d����	 ��glI���uܯ��t���$�����X���r��,����L�4��u3g�kx���Y���57�{%O���@ӵ�W/&�(~���xv{���5<��PH�ۣ���GWA��C�8Ge�k�\C�̂&��v.��L����r�t�*�9<��3T��L��>{)"r	��$((�V9���~�z�P6�|D��菣��/P�12�Hb��T��s;3
�)�Wy]�G*��ٲz�&V��){^��z��g��t��sI��ή��I��V��-29��HN�6Ûq�(,�A���M��)JJր�Z#�H�9ߜ�}�n�IM��y�wc���[���/mWݯ����I����޴���y�vQqN_(i��Z��Y��]�����ۚ�G�D�\f L?Wv&��ɷ!��浉CEƵlW����/��B�:a\��}��D���|S7��0oO�����������B��7���h����V@�xp�;;�Vnۭ3�,--�	�$��:�ٞ�(�ѣ���~q�@�����~��(7�Ǧ?�T��� L�͎%����&;J�F!+�2%��e���LCs��gf�(�a��t�v�^Vgh�����9�MO�:����Pi£��q�m扖�ǳ�ǡ�����S_7�)��l��&r���"z���͆1��de��'5�2������.k�7~�@~7�t����j+5w�x��ߢ��O�lj��!��:eyڧ�7vN&9�ޛ���R����(`q(����D�M��aTk<uT�@�H��U��N�g'[F{@ª.Y���?��QO�Ƭn��gu��3a��r
Ғz�UVB�@��jo�$�l�����#:q,ܡ��+1IM�T��w��sQ�WY�����"䉖��gϤ���ذ�D@q�)�R��)>x�oK��"7$�tR�g㌽�*9�T�̥�����3�����=Ѣ���%K�__J�Go[ۛ���ѻ����N����;濩��sx��U�q�u����o d�d��֦�گ�M�G}eZiBJ�`v�W�*L�|8��\��⨵�������"==]�|���y������"��V�a��_���<��>~{�z%���]�:��%�����}�R�㝂���G�5�������U˴�v��>}J��s~��q����*����[N8����������G������5�ט�����*��š�����_E6��*S֝��8u~�G���#�3�P�y��p5��Ap�8��?Y���
��������z~�2#�"yE�{S}��2�{K�ǲ�������>U�����C�t�D����-a����Ɍ�-�/_>�=L��X-#�ksg���|T�k;L#�ʶ��`����E+2��tt�DO�����(�o
��a}_~�[M�	]��a~" #(��9�s!lޓN��ܝȲ%η-��a撓g2�@���{A4	JP0��r�d�YTՍ�/�����Wd,�o�v��Vzmc#�
�|�츛]П��:����WÏq�7UTx�K�S��?����S��$�I
��@A��h �\Π�!�����?���t�!�A70j���a�w�� ���=�<5�=ts�%Z�ps�wy����F���Z�N�
�^=?�Ӟ��y��m�����Q�iHA�r�<o�q,���7KsZ7&D`5�#]0չ��X;�_X��>��!�TzЋO#O{���d�{�C<w7�1�{*aK;����
�V2p-GY�s~ε��|�f�5Ϙe���=~���&P�ǜ�?�We6�!,W?/C�T�b]�C�h�%*B����-�O}7(#N�i�։�;=�R�ť��hAƀ�J�8����)���4�J�e;�R>�q��?6��)���ӥU0?���,%���O�e)C�.�fE� 4AD���5%�`0�`�=H��P�4F�jҏW���#<??�g��k��1���n"@3O�\3���TPv�hh�7G�2�.��Y�E�`"W�Ö#�'�װ�I�<� ���#?L��5Y�?r��T���u�җ{{�FPi0O�C4fD���ׯ�֟���2/pE�Zu�	-*'��?�
2�VJ߶3��WDA0�U�K5:����c��\���/>��=�a���P�p�)�o?��Xr8>���"Ab��ƾ�_��k��KɃ����N}��o�lm�o=s�`�,���-����L�Z�`��_���Iy��^z÷|9=f9}���8ս�!���a�Z�E&o�7��T�d�W����I������!+8���u
2��?����< VW�g�)��T	��v�פzm��!@U����o��-/@�+��4by��?%<����r��,��N4��jn������P�����~�oi��OA��{����k�k���g$�6�ms���R�#-�I�UZ��۞��=�Lh�B���m��yO=--�3�9�ޡ�Z�c��v��F�=�Y����K	����KBT�y�Ĭi.	D���0ϖqAǭ�g�2~':R�?���T7-�I��D�g	�	�~����m+�W�"�mmvgA���q�6$�Dr��ZA�lj?fE�<�_.	^���u<������
����z�e�Z@�+�mD��#��!u4��`�⒄L��뷁7���7<�,V&����쾇�[N>����l�~�+�urt���U�{�$t��:�ʒ�%�����ր����Jn��`ϰ�e6��w�~�.��pcm�a(���&�t^�_X�0Q��J2�R,f���+M��a��<b0��6wnp�z!ꈣ$#8�]�S��"���8��R���V��!�\�e;??jѻ㡷��=B��I��g�)L�����lYu�ė�Q����C�/!��ȡ��UHŒ�S�WJe�,����:2|Y�-, ����`����^��̞���c<
,�?
�D���g�^�^���w>��T��Oq�9�A���GK&5�i1����-�)��1���� ?w��� ��O�Yjh�0��#Tbej'�ݡ�'��;�|}�uR�l0����dxӵv,Xeraa9��L_�-V�;��m���jIɛ&w;D�/|��q�0�}����P ���[	�7�"W�F�k�-�7�FyW�ΎA.�Bl��ޚ-9P>����H(<�&spӵ��'�bϖ8s���#O�Ќ��Nq�[��O�hW�V"��]�p�p��N:NBd�5�e8���\t���gS�;ю�i�������Be�\��^����=�
�F?�!�9�ۦ�IھO��x!=����d�����M���k.���/q(l(u�hɊ��:'#a��㫎IOt�M��^|lllX��Y�5����Q:x�I?7�d�&����x�/���ux��U��u���\��҇#���qq8�Ӗ��e���G�k��˥��8'*zR�뇒c��}�/��y{��������&Ϲ;�
��y��.�\"�E��7��Kf�й4����2&+0C/�2~���єPB �H�H3����(g��U�![�c�[��M�d��(Zn��s�®�`��q�.�z�N"��&�v��/#
t�rU+�^K]F�o@b���M$���	Y㬀q�\^�N+���\��S+��_7l��`wWg�)�9�+�\f�I?͢�G�=�t�v�dB$���������\777�6s��>-
" �T�5r��}��m���U�������_O�w�5j�英��*�{��i�q�#t��F����8����Mb�I�Yȧz}��K��ѸNO�@-���j�̓M{+z�҅y�a%��Rd�ɤS"O5��t0Q{>(�d?wy����V�Mi��2�C�Ɋ�������v<��J�w�5,E������`��Sw�IF8<�z����`�(0͇}Χ�sf�ϝ�5V��"F��e���F���J�Σ�UJ�@�� �'�$,���[�����Vx��w�=�9	�[�c���CT~/ũ�1���5�3�0%�P���:J(�w{��&j�"��v�����#�L$0R���u���Ojld.��^�Ε���O��&��TU��z�����'�:ϝ����d�o�|�G%��D bV��*������1SOϴ~N��n�p�������-�,[�Jw�6���a��?֯�ă���ɠHp���+2S�XV<$y������FRD���	s��!�HS�"����Ic��<[��ju_Ҽ�b,�m��l��$�W�gk-��S����p����VT�΅ﳧ��ۣM͓��	׫��<I~�Ӎ�z�������Ht��4;7�Tx�S�Œ��3@��.��i����@a``��������-"Ǐ��$�	XS��S�B�߿,֙�TD����,�xTTT���,߳?���������'@ŧ�|�
g�)ڊ"fn�e>�+U�@����Zt���i�	���
��2�>�Z��,�[c5��~����(/����[�6�kƑ�(��2 �����P�5�{���4�����.�XZp��$�Bb!��&E��y��A�1ɗ����1�s>���y+r=�M����O�c�(�F\�P����5vi)���?W���]:5#�_�������d{��@q�#y��J�N��gg��g�EN[l:M�MF�l��ޠ���g/�l���=3gyJ�П2M��`����1X3��6���d�g~�'�,Z��`D"�O��-��J
�5�3�O-�Y�!~�0%��S*�[��o9��O�9��Z����#OO<u|�S�ɨ^L���P���	d��e��Y'1��������XV���IC�m�\�m$�O���SK�!���=!h����i��;'Ȭ��,�=���A` ]����ܡ�s�+d/fޟ�V8��3T��(Z#A��F2ɕ�}��LP��)���jϾ3y��EA4�ÿ!�I|~��}�rX��V4�=��=1Z�>خ�?|��f�f�.��m������Ӏ@�N�.�M7��xAZH56qJ�e��a��MNid�lw~	u�����`�����T5���л��k�И�������_�6< ��p�)�����N{?\o�p�C����� (�o�ě�)I���Qr?V��d1�)kO�qC�>D򥢽]�:`�^�*Xt\'7�2{4r{I�����_[÷�o�#)�#�Rc��!��sl]�Ti�1��_�҄���P�����)����n�sc�|SU����������ܗ�4�	�t�=��"1���m��)�	���l��Q���F?��Fkw���O��O.��pqN�G[O�gm͔���KҪ���Hvσ����Z�Oϩͧ�p~U��_���{��J�Jq2d��~�6��p��@�*���F7�iQ�`ۭA��8[�� r�#Mg4H��@��XѶ>&��>��(�S�ߣ�!(�ku!|��.��k���?�jQ�(�sE��\�]�ׁH��������c("Z���G�G�:q����C��v�����0'p�3kR�LmQy)�u�&}RU�h��)��;X��;2��� �SQa�p�I��l��x���Ã��k��QMM��k�_嶭���r�J>9@�bs�#����n�8��3�xZ���_�>=�����C��Y@���o�\�Ve�X���w65E���}�g@��� K���^�r�\�ZJC~z�O�� -DϞ5@H��K��D�l��\�zX1���&��CG����ƠT��y�޽����{�{���˘������''���>��f������jW�^E�^��˨V�q���,�l�ZM�y��XZZ���
*�
j���c���ݣ(�ds�ztt4�����7��f7X�B�=��h��]k�eo�M��,K��Ǐ���L�|]��0133�ջZ��̙3سgfff��".��ٳ�/i�F%ۇ9SƵk�2���O��(�3g�qN�N�s�ضoߎ��%,,,�ҥK�w�����T*���֭[�s�N�B�lf����)h�q���4C���ܹ�z��z����E\�x̌������:-�8���(�Y}�"�=�!2ײt���2�og(�� ���Y?~�����_<|��J}��F�W�+�2����f�����>f���oI��i!��9�{���"�ipY���������	���s�d��!8���&�A�)~�3/��h��-�f�N,�P�a^3�܀��̏�N]���o�4�}.K�Y�׳��Տ�U��\��n�u>͠2��777�����>������ݻ�W�7C%$I�Y���H!��I��_��������D�·�p}��#_k�~}&��F^����}������m�=�&02�M/x�e��~ԹW���g~�}�/���o��C��D����+��P*M���{��O���i��1��Z�}���ر����������7�[�g�f�9��zx����^�7�ٸ�|w-�� v�����a����Z�M� 6���޿�9ڊ���1���7l��봙~l��4y_�A��ߑ$�����v��ѭr���)���
?��t���?��?�g�<p������o����A��`@�����GSSS۝��)��3�^��0��g�~1�X,n�i}��$x���c�Q������ǯ������2�ES�ibb��U9�@�ݻ�������(S�����Mp�����H�ػD� &"-"Ph�) �Ҹ J�G2�̬ P��-DQ��0H.����:"��RA=�S։�	@���,B*�[f ���v8�Ի��>�vu�F��o���G��ז1�ވ=  |��NXk�*��
�P�I�:�����6#	H� l"�Oi#%Z燄J 3�Ŧ�[!!2V�b�P��Dƈ� B��rf�B�H$![�u��"Rld)�I����zL*�xJ��k���� ���$Pd{�'�Y$��rb��Ɛ1�����K��r�M��dD�0��T��0�a���lL1SpZ/"!bÜ:�ot:SF�<3�|~�K2ݸ[&+6̅_�7:_��^@m")��(�b���2q��`��Doa@K7�d�D4��N&(0C��@��C)��� h�:M�� TJYf�"�Ř6�z$��Dj���B)Cƒe"%�F: e���5�%	��DZ�\E=P�̖�%
z�w�Ek��~�7zI��0zcPD��zgV�:��ט���F�D�fٲm��S[}|���A׉�E��-=���D��d`ź<�@�!�Y1�LzM�"C"J������Y+L$���T�e�$}�D �DqZj#
 �E� J"���A
�b�2E�$ʊ�$�6&k��E�Jk#�Z�Z��*�tq��Y�~E�;���- DQ�,IL�Y$
�c-u���֚����2i����DDʥ�}"
ED($bf H�a��	��Jqgnn��(������9kmh�i��(��ur B�#;:��8���~%t���8ON�(ȋ�    IEND�B`�PK   �x�V��4�� ̻ /   images/7a4be1c8-201b-41f2-b584-263fc50cb409.png 5@ʿ�PNG

   IHDR   �  �   �6.u    IDATxԽ	��Yu�yߚ�r�}����EBb��@		a-�ݞp8��ɡ����glI���'&R��l-F��Q�#�-4��@�M�U�յt-�������~羛�*��7�{��������{��U���}�{_�ԩ����l���4��T=�z�z�V6�fsPI픪�ڨ[�������aj8��<�%C�WYH3��L�9SMG�Ri���f�ުժ3�zs��g+��\�R��&T��ڨҪ���L�Q��Ҩ1���a�T*�7G�Q��^�Z���n%U:ص+5��Qg0u+�v��ەJ�=�>Vz�٫T��`���y&�Ľ?$�Rܫ��`��m�'��*�ʨګ�NoП��*un�~��6�Z���I����Q���0<��})�>}Gejj�z�ʕ��kk�pd�[��[��"��ߵi��Zo�H���N��hX�u��hTvW��.*k��h4����a�oڍ���^T���zke0Z�k�cm���T�w�	t7R�V�T봎z�Z�J���H\���{j �:	ԁE�{��F�{��FN^�Zu�- Vp�Tj5~�|���i��e%p��>>T� �c@�C�*�A�WG�����bP���j�_��{iX�`���~j����x��F��VG�iuu��߹\o�n7���Lw�Ύ��̵F��Ơ=Gc�i�����Jsz�`�U����������Dk�����&g�;v�15�ЀKכ�j���T�����!\[3��i¦������;���t��5V�&��B�2=��15�NM���O�����Tu�h�R�sWj��s�zcNn^�sÁ��)8��mro�a�Z�Vk�Üis�e2�'A@7������N�3��6 �z��[�s����V�z���\�]�f��>~�� s�w�)���uoЫ�S�s2�Z���_c��;����*�Fs؀C4F�zc�6��k4�!�i8Z�v��n�Ќ6���:�X;;Zi_|��}�����/��������XJ�45��ިV���6�٬�F�S�6��f���J�V�;J�]0��h��''����si�֬��>M��Z 3��p��� 5"H��J��̠ޘ�WG3��`��]��<U�զ)�F�:l�氚�Z�GM��`��f��U�pjĔQ{�@=ti�~��&U���`ځ+p�8�
��az͙FO�4K�WKM䓪eҲaeU >I�`�4��z�FY������3�Ju�?\�W{��G��M�f��X{��\��{��'kS��a3��ҠI�6���u�oZ|e���C�����-X�l/[�/Oķ��]S������
�.%ޛ{��Φ�\eX�g#6�A�ҨUa��ҥ�+ w������B�A}Dk�fm4���0�y�c�E�* u�l�0�Z���@�� RL�)��-��n]k�괓J�E�W��C*��_�$�V�V�aT�����h!�9�$�6�j��v��?��� w���?E���fZ�p-�!{y�p��L<��1lT���R��9����r�M�
ʫ�`�HC4�Z����v�ta����w�oH���kmG�ѩv���Yo�#�]IW6��a����� ���F��N6��c��7���ԧfG�ֹ���9+)�흭�;k��;����1�r�G0!8%�Ym4�*���pVEXE �OQ�C���R�	����+��lTk��<��p�f��:,X+��&�n��"������4�w��ۂ`�$�x�^��ʆ�+u80����hyv�mD��0����E�H��/#x�� ;�7��K`�J��^!���br�0��Z�F2�]��z�D�a���0�&[�j����Y$}�[g�MB�K��A/���ty����W�6��W*��0:�����t���:HD34�3���>��O=�p�Ȯ�S�.Y�/��o�#oj�Sn���ߓ�t��P�5��O��޵�C�����J�Ԫ�Ȁ�^���ht��F6�:��4C��e�V��kC�^���:��5��� v������C�3Ih&�;̵�-�A����3Pl	�dɽ�l��M�#�qv7���,��[p��F���r��M��i9�v�E�66�m�#��6Z[[c�Є[2r�;v��]$�t8x�	��
��{�n��h<0^x>͂��0��0�?�Dk���]���Ӡ�{���)�huuuH�Ku�4��~���_�W����'N�Ξ9��c��d��h���2X�IYIk��N�CSb��t����T�I/q�#z��Cw��������_��h��[����la_��;�w�{ߑ�f�A��H���F���:���BlTj �-D�d����RZԨ�F��Ezպ�u�0?P
���f�������.�F��0?j9�J����O�q��Y_�N����ⱚ�:[�;x`v�_�V����0a�ܪ�
H���"+�wSkz:-..�;�#=�� �3V�NT��Fء��I�
�l���1ۆ��W���󎷱?z-����\�k&�����M9 �i��4�X�t��yԅ�M'�5-��6A�477�P#%M��fg[�����]�y��{������p�����7�'����y����f^��[�\<�䯮�;��~�k�O�c�*�s�����X�ô���ܫ;�0�:��۽����qe���X߻w����u��ý{�,>�ܩ����Sw���tfgg�Tp nzj�t{��
7��y�|V�m��F7R��NK�.�Y*k߾}���<� ,*�
�E�"�2�-��faa!���H�A���#�͇\T?�	��r3�*�,4�4��߈�m����І��v�꣙���ph�(à�h�C���7a�1�MY5��u�2� И�������joТ��p������?���Ni��S��m����4]z�4��/_�۰\�4ݬ��w��;��~�׹��gy�	}�������������g����y2�DI��C(+ree%
.����ݯ���}��}�.��f��l���F+k��s(#F0��z����~��=l�رX������,њ�� Y]^Z��߮=�cCr�$ph���6�/--%�.)��f�޽�g�}�fc9x�`ZƟ�p�����ܹsq|�����ŋ^���#G���gϦ={�G��#�M_@{� ��`�]����?���E�f2�tg����>�9#��"�W��vف�-!@��>����"�!:�4^�9Q!�� `HtY�Akz�7M��puZ��ܵ{7��;}����Ϳ�7G?�����t����.S�Fp9�y���0=������>���?����_Fpg`������O?�K���-�kQ8���۲���;�����kp�����9x��={`���3���,�އ~���t(/�o�!�v
Q�"v�ڕ�}�8�ٝ�h����r����4����4`��.����>Ŕ�v6�1�n�׿>=�����o��?w�y*���g�`�xꩧ��wޖ��Xg �ћnJ�^8i7����G�&���ao��栃�V�p��=�W���m� "~|�{�d񮝽�ϲ 7{�tן�0� �\��]��s���}x�]w���;���ѣG;$Q=q��G}t������8��8�����z�M�"�����{ϮԚk}������G��ۯ{]j�^��t�/#�S���z����>�K�.^��馣�Kt�s��j�B=�ēi߁}�[^�����鏮v��ӳ��gN������ޥK�y�w>��cvu�#�IX��r-�V��-�/�|��b��EZi�� 2[���r�95d�L�Yw9�~��J�cCAU������`�28d�-h�X�i^�
�uX��KD�cںf�e*�����z��nܦU@�[.7j�5���6��6��_���Rb��VQ�[nI;w�L�N���߾���<�dT��T?�هv��Ϭf��ި�"�ow������;����=����w_�=\�e����8����깳ggn>zs�Knm%�$h� ·��=��p������1MG�j/_�����n��w r��4	f�&��Hʝ�V���݊ ��qX1���8���V��Vhe�^��[��_��&�h��n(�#���� �n���̣q	�*
���U@l:��4��~,���hܥ���_��w�w�툳 �{y.`6-�ҿv��(6#?>��2/���������7�����������y��O|p�"�yl���B�sp��'Ϟ��sϜ�@$x�?/��{�{~�g���O������瞋nފ��������������nk���c��_������ߊl��y��(�Ĳ�#єQm�)Ǫ&���-�ӿ����b|֘�@ׯ��X!V��a#�b��%����q�Ƹ��Tc:����l@��0W�q�N�\��დ���|�|�y������2L���ް�_c^L˸
Xԇ��(&�7�X��U��1�n���GI�<�.�����;��������MGoZZ\����|������;���LM�^����g�=�tgj��~y��?~ꋏ�N���z�*���E����ﺵ�z�O����B�þ�� �2�I��-o~c�5�������^������G�������w=��*Gsp%g�V���YQ>[9�ґ9u/``um��0[cX+ɊП�N�[�Ƨ�>s��9M�nV;�^@\*���?5�9�y�bi��׼��%�l��ccN�9���ӫ䭼�?Ǒ�e(�3fp�p�����w�$`�����(so7�-Ƽxƻ�g�q@k٨��~��tӠ ��n�ߌ �K��K_:zӡ��˗�����k���	��M�O�����ӎ�����G��󒧯�Uү%�K����;>��_��=���5?7;���G?�?�rכ���W:��M;w.<���C����� �D�$��%�
 $���z(\�
�Yc%Hl�c�������5�m<��e89� 7��U��)r�፿?�m��<����<x�������U^�b|�1�Gc��5u�ž�u7��ny��Ԇ�)�Uw�1�����g���x�
x�*�x7�H+i�/��}~�������2��t�w�qە�;���_�B4`�c�~�4?3��U0'�.V>��z�f��Wi�a�޿���������O��ϷZ�dVpQ��,`�B��H���������������������'��1�{��A[fg�g"�Y��B}bრ�����ejx����������4Rqأ�Bԁ��l��)@�Ӛ&�G蜩�aW�}�j/��a(J 0b���~�j�:[R��<��`��/s�?&��++�V��#��X��/�*%��HK�xU]G��vbJ�Yr�_��~I�r�O&�`0���^�
X��,}�6���dI��(t⦇{$jY�P�u��������0ݬ#�n��}�ˏU>����I~���5�=�w�����~�S��,.�D<�2� #Y����Uf�����[<���kR��o�y_��5����?����(Rn�r@'D����_��Ks�|��;j�c�����7�8�,uX	��% ��X)@�+���\yY�&C�K�Wg���CN�����Q��y�n��a�2��N4O.��l2�
@а�g�cI7�<�7w��	�MIO�(�ʥ��;ؔ�IBoq�9ά,q�D���C�L�8K��w����4������7;m>i��Þ���}�L�g�o����0����'�no����='�y��Lw>����.��_{��������g�x�׈&s����?� p?����++��w�������'�����y�Ϳ�ꠍ��_����ן>}��N���X�`��@�E�簞y�=j<�#����Xw���\}Ϡ7�Z����O�{ En�'�{���`���lq.����'ee�a�'�2>z�e�ў���vYB=��3��%�|�`h@ή���IK&P�wpB1&�L�E.�q1���0�d��g��W�/q|�=�q�:�YTV�ɞX;ELEAU�6p�D���]Y�����S����<����Q�2�W�c5��ݲk��?�t����ľ��o����w���'��?�!&2��(���w}W���~`��٨l�}Ӈ��}�)�i3���2�fP�d������.mԖB�_86�G�XN���/;���P�A���I�ͺ��B"��Ńn���%�|�4�������O�K6��Hs|�'@56 �~Ez����t�LZ@�=��n�_y/�"jDb��-��%������r�x��U�7�ǶE�.��ږ��
�29J����n���t�������߶�4�n�	6�c�(�م{�6p�ʕ<pח����}�o���~�\^^Zt)�\/b�^�-ߜ���w��Fgu�������_��ĉ�Qߔ+s�����11�`ʰ���O��$0� ���GN' �2��
+Ŕ����U�ygu���A�+�4�!E�٘��`�|�?b�*k�
�W���d�1y��q�x��J�Y�J������8X�����U�s�tuf�ysU�����w���iM��l^��0���6��w{��T!�Ὂџ������(��͙Ji-7������|��e���Ѵ!��K˨�w�޷�o���+��4�w�����С���ǿ��}(���]�>�D����8ל�;1�X?����/���3�Tv�H�n)ڕf}Z�GFEۅ-,̏�.���b�5�Ӡ����.J��ݻ\_�ɻ"��H���ߊr�������&k6�Xz�ہ^,��Y7A�����+�Ҏ���ɘu��t���� �"]� ���}.��v�V�˽���b��b�����/å�����"�嵮�&{e񩩼āY��Gx�Ȼ��{.���o;y��#��Ǫ;�8���Ղ�-_<�w���kZ}]�޿��ٛ����g�y���wJ��Ξ;����w������w��?��oy��O5����d�R� KL��<���h��I|�R3��$Ga��G�E���s��n
�r%d`h�J�M�E�֗�5�|en9���qF�!���6�h\d2dp"@� {^��bS7�'�#�JT�{�I"���1�`����C\���O�1���s�{���|�� ���/�mҮ�+~7A�q�W�"��|��޽"<ޭO�C�}|V�)�ehEty���w�yw����ؘ�����g^���zh^�"��lk��YY�y�7_�׾���������F�y�OY�������Cϝ~�飿��qЁ�3R��<�����Rg=D��st��e[����	B%v���<������>�G(�"j����e���d������g7���䃻`�ar#��E~4���@w��2��JQ� d<g0�-�ρ�/��ǱN��8�چln��R���pԜFx��4�^�I��\�&�9�����HW�޻i��՟���=�����{ｕ���ﺀ]����Y�� tn6�'�X\h!|𶩩�S++�U�k�d�k��>-���ɓ3-�E��D�������z��������/}�ᣮah�X���y��Ƅ��
5�ᓐ�� ��V��4VeT1a�G�t;rǜ?���9����@��(���������E�aۭk���b�Կ~l�=��v"g&M8u����4/��bW�ѳ�+�l�ٕ���:rJ��\6�|݆[��tH�+N�����Xp��"���r/f�k����t�_���!(�e/H�ۻ9��eC׉u�]�|W㰔������ df��=����Աc���_S�?u0�8�o>x��W5��D7l���<��{�a�"9�v�J�����0\9��c���W��ڣ���k7�v�.����]2����\h3�ef�AD�W�#L��o��]��sy7�b���m��e�X��\�l3��Ï���h��ޏ�j��6��d͉�[�R�\b��a�n��Xg��Bf2Y3M�`�x�����^N����`Jy�t<G[ۇ�m?湔���Ky6��>dx�    IDAT����O�O�9�g{݋�ڌ×1j���R̱�l��+^�џ�ٟ�\��$�&�1ק����=w���똼��:�����W�ugs�{#�i���TR�Jܷwwj�����4`E��e�Q�VY�In`u0qiy)Ů�̳6�-�6�☉'A� �LC3I��.�6���~��C�IT�n�aC<b����iw�x}~��cr.{1�bm:|���74h<�Įw�ʺ���/������n#f�����8^8.��z�N�Ӣ��nᪧ��t�t+�%��I�W���,�Q�z/����d���nw�L��/]��L�!q�s�������_��_�x��_�rՠ3���?v�-�^�to&��'�����2�|m{�����-Dk�klXJ�����+��8nip�����T� /�AN/Q���bO��s+���*��ƈ�5��P9�w��9̤=��dw�KT/�-�4�	�{����i�VByqe���p�W�yg��W��{Y�Ȋ76$�̬�(*o
Q%��Μ��7�]YM��N�>�����p:��P��v����ŝ�m�̯9t֞V~_�g�,��4�[�b���~��~f�~|.�x��~�]���2:{��`���`��UR�w���f��;�>y�q������c�f��?���7��9��G�E�<7�����'��X�����o��'�!���*k�i �6��c3QM ����	�D��A|OЍ�F�FL��_؃�,=!/�z��	b0�?f���d��U��\N�;���r�V��_H?��ߛ~�'�}oL��c���z���;̬�7�k�c-Hħƀ�=������ ڣ������}��!�O1x2=�!��ɁhЇ2+��eؽ��$�^�[�z�Aclo����x��ڞ����a}��ƫ�gY]Ӯ��/}	���i�'�|<T�kk����;23?�.����<\����]o֏*7�(�����G�{�P�͝;{nJ���-��#[��V�пkC�ɀ�Z�����G� ��8஀1TS������?�j"B�����B�i)\<89y��D�=s�R�;?�w�;�y���׼P#J�Y�ȅĤ{lx޽�^0s�e�+�9�!�� ����g��w����w��~��>Ė�+�j6����l��W��(�n�4/��!�F�I��<��:�=���%�k�Z��-'Wl{�G�?���c?�c��[oM��ǂ���vгէ�կf���3�v^Y]�ET����l����uZ��ڕ��Ȓ"c��F�u��r@��a(Q�~՝�0�;�t�W�� 0:jE���c<2���8gH#��Dp�<K���A8�$�O����Jٻkw�����t{#�G~$���X^�H+4R1M�⍃C�:K	f)o�%Ͻ�3"�u��"����^��q���tӾ�閃G�/$;�u�?'��^B�xH(�$G�Ř�k�'���k�y1�M�1��{2~�帓F;/M���cq/~��]	�B`��Jw��#I���ߟ~�~ ����+1�T{��T����g������6�iHC��NW�?ɔg3r<Qj��խ��͹ʩv?�yӖ��% h�W#s�1]"��ݳ����,U��W�^���{L�D0DD�=B7q}6G�ʂ{�?�?�~��~*zOv�ݧ�v +�LM�R��@����Js	��"�2�6lv�Μ���"+�s�3gӷ����w���c���
�|N�=݆��5.e�T���z��I0Y�k�O{��)�-���Hw2|<�G�>���/�|�L��Qc&�����Z�݀����/~1@���iP�_`�Zm���5��=!ou&� �W�;v�sG����÷m�3���򣜫�&EZlp��^F+�xg3� ���\B����! �HA��n��wWgi���Nd�96�J%�F,s%=t�6��\�cu"�I?��ޟ~��ޛ��?�����/_f��q�+�zZ\��a���B�O�G�xfc3皱�� 8�"��9!:��Q�NU@�8~2���#���ߖV�	.^^IQ�'ϞN�◝bI�;z�Ln��c�y/d<���=�ԡ�6(��*NbB�����qz"bO�����u`Ᾱ���tB\���w"cP�d��;�U�+��w>Bw�"ꓞ�Cb6����=�G�%�%r�jS��^P|� u���<�ݿ'�20�ڷ� ���$�z���` ��\S���[V���o�;j����ڿH���:�I�R�ܙ]��}+�פ���yw��Jq$.�U;�ڈ
;w��xn֚�s�A�_~�{g��U�6�)I�R�ڳsGZ�t�6��e�2���X��(��UQ������:*�U� �� ��,�an�R�f{˂�m�4���������|:�z�5&�R����r[Ȣrw��L�������	Ĵ%Mt���k�->mi5IG���V�H�Bs�͠��`�r��d\���	46ƥ1L�d4e�=�=��=�Ju�s��&���m�~���PGG���y�Ec��f�v�S
�I 춞3���eoȫM�G�$V�&��zZW��9U�l'�G��V��8 �ҕ����X����t�]w�!.'\z���1���HZ,ɽ�]��}�|ZcAm�6;]��dznW�8B}�͙M1E��M
�9T;fgL���F+����3�G�T������ԌϞ9�����Jg�.�U�p��.���E��Z��^��T��aB=WU҈H6���Y�A�U����M�n�=ד�'S(�W0@j�$�����'�o���GJ�(Ø�n�5|��a}�4iykLt��aG���I�Q�jm�ڵn�y���w��<qb�I�>0�=��9s�|�BX�R��,h,dl�3���E��eL��;�
�L����g�� -&�bU'�._:����7�����I���� �9��tGD�H���u���@�����_XS/�����`F$k�����W�퍛I��`�TnL�s�q�Ip�*�g��K�2х�2��uy��w��">�ܩ�O2=�����w�5�K��w�#��W8����$"4�<�cj!��wa�a��H�B��,�|�n��:-�wK_��R�M����\��/�3�-v�UZ�=D4p�h�Vf.���Vޑ����y���>��K�R~������!���tkz�aW��Pg����=��gb���(�<o~b0�����j�R�%�<��X���D*B���kz�h���5�񹲲�J����p�}1Y�L��ƨ�Ђ �yuWN�J��Ҁ��2;��h:jk�����BL�BC�1�x=��"��R�yP�i�Gn�����?�D:�[ED��Ag���e1�-1�D$ٍ۱W�*��N�G���O=\���Sy�M�u�政PQJ�lț��!�Rli�I �n�+\�pk���1Lwm=:�)��T� ;��~�?��������Z�-�:�;��z�'�2C�G�՞��*`ɉ^����MfGjC���AFs3��啥E�I�:��p�(�8�n��c��[�i1�.s��	���Y�m���]{�&�𨁟�'�8�y���3'�4@�Xe��3�	Q{p�S� ���p���rڀc;Pu�X���Ȼ튬��iT�jGPq�/�_�#}B���A��H��M��80���{<A�u ,�bn@���6��t+{뷥{�}]�(�?{�f7���W�*���X׫�0��b�i|[�վ�Rҭ�W�:��\W����D�J�"�M������K��p�˭����^6��uc����/|�~���[���Y{��z�F7?����}3d�A
Q��N��~&���	Q�0�K\>oAo\�lY���� ���� p���q;vK����u>~6��}�8_h�S�{��kp͓�}9�/�O�����Ѭ4��S,5��0�߿l����"�Q��C�'r���54B�;������!_ I����J#08�>��	����[̊�h;쭧=��|���6�z�p�̗K�?��\&����'�oV֖kKK7c��xs&cis�r��������f��>�V��h�]x��lH9��0d4�g������jL1R�J.$sבu��n���+`s��a�x��~��ʕ��F|pe����& �#�k��HX�( Vރh�W��W�L�+��ь镟����M˖�@<+����-oyK�G?���Y��h0BW>�\�s/q~�n&d�?�h���Ӊ�T'�,��ڼ�m�В�9�ީq�lҩ���
RW�y<G��$.E�S��&NդV��ĭ1S�R����O�?�h|���f9.Ã��hI8c�m�i7~j����sHP4I�u40�� �T��Jm�"����(�zy7/ l�.�:�9�W4�q�e+�\���S��ǖ�]{����)y�.>���������ǉ�����upnN���8g���ݜ�\�6��w٧�n�L[����֮�*;�LI{Av�w"�,��rU��6n������/��ϥ{�]/,q$�M)k<��G�F����s���=��� j����i��5w9��	`��\UY�� 22 gZ+��(|X&]D>_ر��E�@�Z�/rT������6��a�3����~�i�H�k⦶D �)�f}*��*��`2�f6�~������v� �RS�C�y�x�\C�vG#}��u��*���>y�Y���2)�j|πͽ�n��g�Xb❚��d!DF���j���l���zm��޽/����p89����B4S��� �%[���}�p�K*-��׮�+�˰7/�{m7�I�����ݖ��?��t�+_��,���C$oʦ;��,8O<�x:�g��9 �gQ���"(׈���@jED��8���LZ�f)�x�7'��a�e_h@�sH�N���K����N���,	�R>������"+�X�AW^������&J����Pi��/|�ߗd"��R��_��y�nU�t� o�{a�����T"_姸��r��^6�F�g��Y�g����n�\e��:S���1���Tk��Ũ�77̹I4F>N�68T�c����f�hip�b��d��f�6	q�FX���X�r	�sӄ�$����3Ǖ��>7�/?��;����'�����4`���g>��t��ϥ#�ȧ \zp� �8]8��r�=��gʕ��I''@�4S�3i�!�Ѐ�j3<yG�H���x�w��~=f�؁���j��`�\@eAN���~6q-M�M��V���6�r���}u,�������S'��+i`K�]���+!��%<����h�lD�VSh�s�؇�Q,�N�r{����f���
'��	����c6s�����ZҎ7A�r�oݪ��O��i�I��������	�L�=E�F͹p���%�����N`1&�x/�;
[(6�/a����7���W[;���E���ۿN����L�?���S��B.?��G����t�-��>��5��2��2mL% ��Tī�Ь�����9����W���'Ʋv��!��@`��9dcW����s|�δ�N#
]^B� �X�iL��-∹�>@����w���ѵ/�:s�1��-]F��F�~�s�Y/=|�Lڳ{1-!�HJ���1����y��VM�4�7	�C�E�V$�ա��2�<gcrح:,75'��lk�,�|�Dw��k���-Y���͎z����ʿ���d�hV���lo���+�-�o�/��F�c. �Lɸ">?V��3C�iL�#�m@?��M?�C�M�;L��Չ����i�w�s�O����i��*�r����. c�%��D�wbG�yԡ�"�X.��+1o ��/���j���������i���YH�j4�MT���Sس��R�B1��Qp�<1p��Qıspp�z	�3�����T��5*D,�^f�ٻ��c�_����Ef3�\[?g�P�c�1�1C�\��ľ��۲��M�1L~.�.I4�N��l��ڵ1E<5�ůq��G����{`�C؞�tN+���$εK1��K� ��(���k��ߟE\q��#�b6[,��b_�`���Z��7i��~�p�U\z�ь���Mm�N�;HSgܡ�����N����ʙ3�>=Bg�d̀uʳ�q�i	hMɓ���zS�U�,����q�v��k��^͛�tz����QE>�.�.l��ľ�H3`Q�"��*.�Jaa�M��ʙ�
Ո��t�|�5�m��ťt������ߙ�Yܛ�<r�5�q/4Y�I�����?�5��+3�l������L��Y23a�~\�>��\dKT�M#���ڨ����67Ĺ�҉v8� �����n���Y->��(��>s��-Ԥ)n4>�4�� ����0�%���~>�t�p���^���Tn����G�U{?Y���-��3[F��"('W�l?��ט�9���rN���s�1p�B�p��` �<i95�;��B�^j�A����q���!�Uq(��^e]>��i��KT��� Xڅ�S�|��o8v';�6��J��%�|��T6�7��,�VM��\�d�����~� >ק���a\�<WX�Ӵħ�/��m���eE�YcsL�5���������?7���m�Enؽ�~5��8�&" ��J��M.�*2lzɅ��AhʩT�7���F�NNeoFăa�f�n�@�'���P�~:��fn{晧ө��J�3s���I��#���Zѥ"��GT�@�2�������L�Ϧ�Y�vd�M
G^qs�߽��*��U�ˈY�d b�3�ӽŠ�M�tÔ8�y�&\U]e���j�(0vP8B���&~^�� ���ͺL���W��N���/=��	��ӈ6�g{/�Z�����b��t/��=ב�����rz�����l�+zD���
Ӳ�S�]���W���b��;�!c�{>�__k�EEO/W�\U\2kf�e>A8V���2��(ﮃƖ��N����*L�G��7����w����ҿ���v��B��b" �Z����@����'���� ��}�tϤ���d��3rx�o�L�z��f߽L�����=%ki�u�s�u������v���3�P��5�c5~�͌'J�@���%�p)�K>�<b���P�9�P��O���#�D,�4n��Aj��F���M�N ;s<�lV�[�I�?��t.�L�-�l��w�˜��ft�0�
=H��g��!����uFP��ɍ���a�Ϟ%4Y�ųV��?��`Q�GYۺ6�b���qbt"�"T(�.̥%���Oͽi	w���`���;���N��i���S�=Ϻ�`,Pf��:O>�>	t߷9��'*����W/z����7|����A'gg�d3L�4���~�QA~�T5��hE�Z�l�K�fĢ����@� NTI�/F\\:#W�n#[��3��ʠ�"{�wltJ���U���Ï�8�3����U�i
=:/َE�tZ�U ����
����N�O���34�@q�=ߔ�L�����ʈ�#l�� {'��C�S��̩��t6O�6��y�V������.PK�J��ٲ˸���|���.N��=}�u�d��"�<C8��Z��&s-��[\Yq�w�x0{�6<�Z�@�]�f�f��]Fk��
��	]�m�]n�z��1�,w������OR9p*����,�b� o0�|���=�;p�.�dЦ!8�)Q��)6 L���C�|>b�h*��;�B7:�1cRn�������\��o�����E>S:m5/gS��
m��(�zQ��I״����u�������\���KM��Px�
ǐ��S�<�q�ƫ���
�����q��C��;��bV���4v{F��R��5X�jg=�+���."����L��r�}�X�\e���n��]cʸK�]$5@��š��jYu7Y���R�R�r/��%�f�m�>�+W ���=�r���MG�
��	4'J�\��~ .@ѿkܨ�    IDAT���i/����f��mqn	SM'0<Mν0�p��#��=ߛ���J���Ui{Ӳ���XcA7�E��Efo3�ƅ�U�+����_ ~�����ao�r~�rN��ڕI�2@��8��q��q]9]YhTl,�o~�I)z�3�E_d���wߓ承Όh����d<�-딾�6���178���D4r�|�-��U���<b	{�5�nK�N��l޽̓v�b����5+��^�ܨX�]-��a�[e�-	�ƭ��~/*���[�R���{)p���_q+���XKN����^�'���o���1��0�OV>��͌��O=�N��ob���$)���h&_������U�jw��n��hɩ����+�Nm@���3�ɘ��)�A��6VH��^f�+õ]�!'W���$�w�1�֘K#���2�&�!wg.�o�3po��Y�z��'�����xi~��4˦��L�_�1`><��^{���矤�6~~�K���.�BN�L˘��xъ�d� �ԅ��f��8���+������ɺ7��.ǖSkWw�;��6���Ԗ��D��~C��ر���#id#�6�9Y{N�'��{K&M�dz �1�^�5ig/My.�aIr��؁\iW�!�����RbwP��S&����g�MSI~�#��QA��=!��q�������m�#P$N�Lm(������Sl�=�� ���Ɣ;u� �ˠ���U��C�W~ﱟ��������ܝ�e�<�P�-]A Y���"��&�ɷP+���;M!&bG���=�qc?P��2a48^x�D�P�o���txa=jG��a�̆�T���sQ��2`�N�q��y���K�}�2��W��O^�_	��������ۚ��wم������8�?�����(�ҋ�=7_f����R��B������l���}�oy�C��v}���l���O���#S.�f�?�m�e���4�� �%����If�����ʼ��Mk~G�^D�/�ٟ��>�.��\�*�ԔAϔj�n�@�*�#E��T�2wpb9�y֓�+8�j�dE�X.�xY�(�BKa�pC���Zk%��(�Lr:ζ�]�p�=;XW���f�:y���M	���8h\j8�7i/�=f�x�fo��8�sWUɻ&��{�����.#�\۸��4�����)�L��h�֎��Zn�!p�l�'S7
�Ի��:�9v��NrҘQ��/�.s�ܽ��hW�OƱ��mGV�'4�wя��w�}�S]�+ru��C=�?��8B͡�jЭ:(� �xT�~��$�3�. ���qR��1f8�!ו��d4ʣlh�T��+L�;Hko��i8#���j��ĲE%�3�̣?�%� �q�+ ��0į�t��v���� O�K\} ����9�P�^��Vqe'�ܱ�{�|��dH˝E�d҃6���U�d}�z�S�c�N�{�a�W]w�uJ\%�r�wq3�Ԟj��y���/�����ùy����t�����z��*�n�*א�Z�Gf�D�ϚRHߣ°�^�����8TMł|
mcz���S�����T
bXy:��3ibՐU��7���չ��9�6N�i�Z���No�����t��'B���n����y�yF�����}w��	�yf��W�bBrC��(�o6\Z�'�hq����co�p��+󦆈(�D6 O��!�=#���{���m>�t�Y��(���i�<�� NZ�,���A�;�O���[��R��;9n��Wȡv�G�bL��u��8}�2{_�TH�D@�t�*��ue�Pyө�h�X����(N�8����yAQ)LT~T[k�*�gk���q2��O���3������[n��@�XR�Î2�X
y�O?�R.@8��E�-��AbG��C���x���)v��%���W�F�md� ���K�|�
p�B8��8�3i�r��q�J�ҋ���#�4��Q����[����Z�ӈ�x����Mhd��?����+���0�<ɦ�U����(�)���:$��ȏ�Q����u�яW�� ���=�O�(G��+J\���ɸ��H�qVj=�zis]�
~��۴V�YJ�ϨߺbH9>���_MJAlW7���3��~�Ζ�&�.ݾǃjv�)`�~�Lz�G�h�w坲���A��KP� we���ݜvt�7����<��vz򋏲����&q�%�6��sPF�!V�8v��3셸���+��	d��gG��R�B�ɻ���+U��
�bo|qR-���v�� ::ɶ� �Nt��=�$���%ݼ�u�g�2~�C�׏��&M	/(5Qd�1mC�~z%���{�k#�VIbh��p��:f+��x��f�Ih�A8�'�9
2x����������)v����ɰ�LBU��_f�ȑ���E'\ �����I�����,ge1]n�*�Q@T �qHe�D�ͺNd��G�Y��H5MsN�i��C���ś��k�J(rDu�+;Fz�l/�&x�[���?�w��4��,4 E����e{�6M���8{�	T�zu�*�m�r�+jq����|������E�j�L"�@�ٴK}�Qy�*�͌l=�>�g����WBL��^Ϯ����r�R�L�,%�W�o܂
}>E^�.7`?���[\!BI�d�B�����ݏv��a���h��]������7��8�	9��+������	&Ťj75%�H���{A�I�@���7Ϡ]`�b�"�hQņ6�M�R�Fg���@�b�������`	-X�["M$8�)�[`Ƞ7�2��F%�n�c�θQ����A"�� �Ac�}��ZCd��|���сY^��!�A�n� ��]7�� ���36Je�h6����z+�.T
wk_��ʢO��('i��1�s(�)>Ðf]�y=s��~�=;��9	1��X�&�٬�<f�
��@)�ϥ �7�cEL\ž�_�o�n�������@A���'O�8-�t��2�3s�>�E�4M]�i���Y���M�z��SMO>�t�Ϟ>�P�f"��RY���x���&rӍro1��\�F'MN;7� ֍�5ʝ��"Ϥ3�ڦ'���lM�ȹ�(u$��l��=��g��L�jLu�'�vլ��x���I�����{ɧ�r?��8���S�;�u2J���<�q]�7��b�t���H�'�+�fƶ�k&	2��]��-�𺖮��4ۤ�=����Τ�#�xq�;֕o��x�=�-�w����dAg��\�[�qڻ_��G�\.�'=���9��p`��,����w��`����+�W�.Wu@�ϨP<x�X�b��B?�!BO�#��QN�J����G?��~MŸE�Cq��&��D�2��L�g.��g�2׭��ix��q��ٸ�Ճy�e�b&ӑQ���ʻ���&o�,��4��-�]�����s�K&<��%�.I���xŋ�����B���|-w��3y�21z�Ç�~���1 ���c��r3Ƶ_8��L�Å��L�Z`X�r)�LS������t��[�Y��i�W��C�"F�(s �J�y0�B�(�؟v��i��'hS�Z�O2������[���mc�!D1�SS|q�w?N�#Q����3��iq	h/M��~J����h���̻v���8�S���W~j�u��y�Q��_�l��K�����{��vB��$K���Ff\BJ��Ѭ�v����K��5o����X�IfA�0��|��f����"m�n�Ҡ��[�J���p�&�$�Y7=��
ʪ��q�XQA�l��G^%)��>�-v쬥�_z(�X��]:��z�xUM�渂4�p!�#�嬔��6Ċ�A�jZ�4Uo�Y�O�sY6�:rw��=hå!����ʹ����@��>c׃��6�lE��{���:*�
c�a�^�	�9D��ǭ��_�Xb��K��]��3��Lk�x��@{JFLs��}��ֱ�ԛϹ�sc-X�R�/�R��N�?�u+N<��g�&r<�vֹ�mϼlK^�����N�WBc�w�62j�hJ�-���\���G~���}ҭ<O��l�eiL��FQ��4kN8/�]��1�c#�1�/?O��t���i��<j\�R�h2�v'+ *�4K�@U�+ؼ������!�G��4J��g�n�z�q��R��U��v�<>?���+V���9�Uęqן4*�+qz/v�^�,�O�'�M>?��G��%.�Q�CQ�Q��/�3�/�z�t�}�;uO9�6�ġ<%�ϓD(�*�(�X���(�fl���e}�\�V�����g%�� ��p6.�C�W���
�\H{�:6���MԂb���v���"�U�g��B
7�3����@�d�GZH !y����R�Є8�2���3%�!�O�9->��`�N��<�Xā��YW����yv�	�0׵�W)W�Ǧ=R�Z�-��{�W�y/n>;�_�.�O���ne$rx&�#/�!=��I#J�fs��4�Z�&:mz�8*p�E=��@�%��^�}�c������]����ɾ��5����D�I, ��#8 T�[��\2�C��U#P �Z�k/ZR40eU��h��2ĄqE(�X���E<%�F_��x�x�L�d�Ы���d�S��]���n�vW�C��(��9zzo��~Eg�����2n����~�5�=�~J~���v֭��g�d�ʵ��Թ�'*m2��g9��lj��Y�s�(5�?���E��yL�YcQS
��@P��F,�o�9��x�	�C9�D`XeȲVqAbL�.�<P���]�'D��j���,� ��͑����R]d
~N�8qt�o�T�m��z�9�oEY���%��(�"å⧔�<���W�6�I��T���\�Phf�qEx~�mO�/h.s	�t�Q�{��'Aܹ��Uc�d��uoyʏƭ[��0���I�4��F����e�kv�<����S�7�ڼRn,C��	�~KW:�S{dC(��t"%�T��&ʜ�qb_�Ѹ�LF�+���h�o� �#2f����rq3���+��	ϓ�RI�ʗn�s;Si�jI���q��(�nu�+��X"1'�c�]��EOd��7��A��`l��Y������]��w��E��2/�[�?y��ڦ�ơ�v��1"�q�tӽ�*<��n"N�1;E-�{�߲K75.�r�jQ?����f6B\RtAl1я�c4a��U)��%���տQV%\�7o�\��f�����c3�R�=3��Ʋ��2fHp���)�'��䙕XfH���R���R
:i��/�p�$������6�-Q)V�1&�D�'��g��j>W��K��	���p\p�yw٨������o�ek�vW�ɉ��+���p�r9�x4K^�Lp+�N��`΍"�&�"�d�uW����ރ��1��z�HO����!��qk�	c�^I�k�盎Jw�~�xL�'�[��l���0�r/>�~��-��>J|宨��l����E�my�#g�q,_B���͡�zy&q.^�Wa���5qN��۵#y2�y(��n�BD�����$����s&^8dhS�Icr_-����0���?z0*P��&�<��6tYk|�����qؕ:�r��KC�S֨�膛���>��<ΨQI�B��ڱ��S��l �4��%F���b�Ʃl,��g��J�n����2ZO���h,�߸������r��.u�����LXIE�F�S�(�n�n���a&�e:y|�{ae��Ϙ����ɸ8�v�<;׵��Fݵ|\���1�v�og�x�-�x�s҄;)�ٳ'�c�� pe��1�Uc��Ӕ�o'�����f� ���`[��J	VTLTkT�r���k˱8^l�{�c\�]N��ӓé9�r�J�AZY��G��e�h��Rc�wcn�*����Ԃ9-t�Ư~z@���v���;�?Շ�P������B�E�z�7�(��vY6��Ǹ��W�uP��H�OmH��6Fp��H����#=�W�����L3�DC�ԏ��|E��3	҉�!��`����ə�তY֠h��ˈL�׆ g�i��ш�ǽ������2"ש_0s��
�\��K�� aͤ�)�;���`���@.v�U����Le�sL���@	剪����̠����$;P�Ո�Y�sx|� ���\�P�� p�X"J�h������i������8g���y��L�7���J�of)0DY�Cɿ�&i1pl K�B�w�!�(�b�8C�i��pDilҧ����|����>f68�\��p�ݒw��c�����9iv��RZa��	m<���G��,�-
P���^;�K1�/X'�v%���Y{3i7N�d\bi��h4�hM���ű��:�x &m��+�p{�neuu%�bJ>����	��Fؖ��Z/��LU?�g�}\�ؗ����m�!�nN�>w߁�|��I
�u��:��YGD`됭R4��д�]���SE��w��;�O�[P�p��nK~��}��1΄N����qܑ��,��	=6b�x��g!���UQ��'	�f̥3��⢖���\���a�aXXa\�H]�A��p^փGħ_�/�(�s�l�L^A���.^����RA;Mq�~�X3!�ذc�!�)X��?�ȱ�<F�+�̤�g���p���V�/�$� K���终%C�s賶#87*�ؕI3 '�[]O������I0�]�+[���C������G�����x���_F"�
� �0c�����G���Blh;��-� qҳ���=�����5�N��'��ES�`ײ�c�{�A^�:=�B|\�5�S�0���p�&��|:\�v!�s�3����)��p6erS�1�H� ġ��nQf�!)�`l��z��(�,�xx|��S�߯/(R�µ�XS6�n!������A����+~J��x,"�'��/��ӂ#���}��K�G}.G�H�գ}87;�)�{ �
rni��`8����%��g�-��z��3L�|���a��sQ�\�xMO�H��̉�-��^����'3���p�9 %7�3�pSzF��4z�~�<�A�nPX9u&��.��l`��j�@ˣx�g��вxn���ß"_�>*�Ԇ��C|�Sк����Qoƣ(1C|��u�)�'����7@������Lm��1��8��J��K�r�i`jn6�O&$Ի�i+�L@�,n�v��i:�& �d�{�cm��x˞����e?9�����g�A�Ϻ�@BQ3 �/������p�h��c�w������")��绗 ���,8�-
o׶�X`�)���Y��׏�������A0h2��!���Y�	��� ۅG~�`�])}�y�*f�#4���8��1d� .#j���\�p� Gu#&8yU#�D�i��DB�H��� �
j9���*���y,��	�d��%�=ӌؑ@��ir��5�=K4�.�q�����c��F�#����{D��+E��ORc����3��o�K}�z`��`�4��LS�h�[��؟��s�My@Qư��g�[i�c��٨���e���$uɚ�{8jJ����%z�Bܒ�R3�cEX +�g)�	'󿆑c�0� sx�k)g�S��$՛o:���
�?�#~����Ө�:��z���tQ��N�ʋ�o�y�ݐ{Q�O%|(��c��` �,�5N�m*�S�~y,����3��Ď�U������~�2��թ}t�Iy�U��#��q�3;�1c��^�g� rA?����� ��0?��'B��':&�G�6kh�t�0��]f���$�H>����q���"�[v���u�U=��&�e����˰d�A;�牯>�2�vݥ%����"��}Sv�t_�OM�%�L���'K�5��w+�L^�X�r��ͻ��n~\���J�RQEbԘ�ڷo_�}���@�.��AX������d��;wO�m��]�\C$�4�s���'RJ�,�*-���=~+�ˏ>��'��)�Ӟ�F�6by	}8eS5����9�(�    IDATw�3=�g��&�Hs���<��_����3ir
GV���7N��UN/ӿ�C��(��ʹK^J����[�_{�7�����n	v
�W�c�m�9�_�hO3�6jN���#2!�q	�`��+b�@.��O"L3o[�B�)���R�Cę������#�.���^@>t�P�g��X���ඞ�z�Uw���>�X���'��/��Q�H�/��a0�"�n�A�z�mX~?�md����yn�K�e�93{����_��:�uv��=�:gyZpw����؞ECq�˜'q�)����g{����ۡ	�Z�GS��:�I:ƹ�p��F'�e���i�o�_|��#t�-NЪRF�J*i�g������J�/�I/��-��ͷ�~,���y0B ��C޶��+�(^Z�>��Y�ʍԼZ��ze���jYT��$��4�����9
O�̈P�s�Y�sC�~��^�P��ٻ�@����Tf!l��R6��@�ZF�P��R��w�h��IS8�r���zF࣏>�n~ű���*i��c-Lϡ��0Ts{w�[o�5�<�t�G�n�A��g��t��G:��G�t�a$�XDðB��k '8��j9 7�7ה�ʳ�=�S���F��i�:�*c�4͢,�Că��Q�Vz�b� �F�=��ic�*^cORz�V=U���t����;�ǂ$ft9��A����Ȅ�~�a�'�H$) �?�j����r��ز͜����Z�-�\��S���������W�rD�K������;W,�hz���+�LX:U�Uo1��P�̖�����{d��ƻ��2�	O7�lt�����Ox����/����BT,q�T��c޹/���4�§�l8���НU�!~bC�+�j��˙U�
��a p��/�l���,W�ָ�+� 	��PM���Xbu��&�'�gt�ɱ�VΖ���xl3����"�q-��	&��l���uΰ{�cS�Q��똿�Ӿ���F~��Qz��7���z�g� [���sg�rZ.e�.�Y���N{	 ��)륷��>s�Ro%�ڗ��]�^�n�z�X��b�b20�ʄ�E�����z�O=�A�!s�9����pfpi�@�Հ�� r�$7R����R
�]�܅�Q��Ʈ��%pa?w�8��[_�^`}����St�뜫� ����S�Z��=��9k������V�!%%�Fqj�-_�����p:}�SL߻@}�]�b��{�Zŝ��nڵ��q�B^']Lp�@�h˕,p�q�N�t�dތ��l �F�jԸ˲��1`<N��Q[.ӀOP�5��(*M�Dx���#�O�n�o�W�iO�U�K}��2h����F&�FFw�C-��u�������;�b���9�u�1`0��L��>�	�(�d�{y��h{hݳ����y~�zS�zU��sW�����HcG5& *��W���b\K$�J4ѨK"*�(��Lڤ����z��_U�y���y���߹߻��۩s��;��>��ϔ6�����d�}
���H���A��>�����X��`�Z���_D�}�fX�dr��#�0���+}���"�2H�hL�K���Y�u,��!F��ƕ����h@�_�}P'���|GrV�K�}/����:c��r�" ?OZ�Y�BP���R����o��%�o>�!���Am�� /}��.�ZX�ݺ;�a��G,����h�*>��(6�+;#/mCf���F�]��9X�!u�0�ԃf�*�W�];@��s8�B�-�����'���L��P<� ��my��`�[�Y���m%U��.�\ i>�я�?�]"��$劣㉇���'��/{�|�?}�����*�ts*u�G��&�,�`25��s�	�GZ^M'Ւ�P/�Yw�<n���*3x�3HK�GX rP��fGل���byy�C�� �>__��`���Y� �#dx�0�ut�����:�A����*Y!�{�=Y�ztB��]�=|�X���B�xɅ/��0ccՃp'K�z����k�{�A���6ôv�i�a�̕Z�T)�Ç���¾(�[^�)����ujXǛ�!
���������~�BwM�n�Z7%/�ҕ��a����,��Gx)I�J0֘�XF؇}�)�� �#�],q�`_J�D�ᒼ�|���W���8��4��Y||@�m��C+�E^�6Y���p����S �"�]�Jl�0�-\�E��>�7r��<[����;9B9]��CHc�apsQ�IsS�.�&�vz���b�;��D_�Ǿt�
�ȭ��b��TG�(jt�� ��.�ϰ����/�y�+b2msQ;����v�|���>����n�Y�c{e8ͪ�g��W�~�io�%"�+4��E�r��N�+��E��? �����ijހg�Cꬨ��TY)UM��?�2h�0�n:�q��4���y�9ܘh"6
�1���d�f؞:r��~�W��ѣe�]ւI�����#���Tkܫ}�I�AX�X�!��l��r]t��6�:�r�ny���e�r�0Q� �u��c�2}�f����W�z{RF�_���+3B� �HV��L"�sZ#;�|��~���kR��W_8�pǟ���뽇���,���BG�'�!���m�L8�˛Ij�ݷ;e�$��.پ�U���m��n�*èˢy��:���y�j�;��rOL,#�������B'E�Rڦqn��%�fa�w ���'�Z\��u�0�9yUW�n�2������]��q �j�`Ec��9]�X@�`�v����2��K׮č��<����U�e/׼ʅ��D�ʮ��]�����GG�����T���ػ���s��6oMn�@�7�P�z�*����k���W�3m�.��2:�$�g�}�����~qF	e�hl��X�P���Ġ��/�s�/"���D9}�s���˕�&�Z`Ak�Nw���^��˰4�,:���eǰ��َ������[{"�f���1�Ș��햺a3\�t�e/Mϸ�{#�!�{��u�|��ĸ]��2�;�}!�i!-���n@d����S/j�(i��w+�*+�~	�t�-�i�c8'���+����z���������c1���y"��qx�cg�+�Ǐr�p9y�ly���r���-.���$���π�Wi��R�5ʗ��א
�xuӮ<����s���4�2�]6�F���R��$�ӷa[�i�}�ߦ $�q`hHYt��*^<�]�f����}�K�Ɠ4����{�9ɾ�C�+tD�ܸL���!��Nr�䅛��o��r�:�� /��'��u�E=| �Q�w�{Ͷ]J�tT"h�n?u��?_֖lb����6_Z\��`����B�����l�fN��(�Q{�!W��mv��j�6^kP-�Ɛ��.����;	ri�g~�g���
��\ElJ桪��{��-�'�)w�yʚ�j˳/�o� �i�C�<Z.s����\b_ƥk�� 4&����sM����:��n�{��D�94�����:>H3���Ç�}hk��壑ր��,��$T�����0�ց(�v%S/�J�������3L����۵n��H�Ν+k�9�|��r����CW��Y��2} ����*�!U��z"�f�9�k��j�gx��z��ba�n}��s��񡺵:��g_�=>�Pg8��̛iv�-x�����`٣���ej+4XƬ�i�q��g�D���K��+E_��̓��0�[�E� ��������̙{}8��a�����s����9��.g����Ʒ<2����(\at�gEs���@4�i)��?^�����;0`yُ�7��Ȯ�� �pc"�������8Q����U/�߀�wQ&���o��j��W��u�g1Ǐ-��=��mwvЁ��n�C?x�L�f�9&������_�^˪�����<���P7/�6����	�k�l����@K����K�C�/�7�YgU�1=�V}y����Vw�[���˰�я��S=��Ą�`T�E�N�V[Ѭ�z�Z{N=û_�m�����ۋ|�k��B�?��r(�JL�\)�}��p^��Ξ.�O�D��U�9ͫ^G�3y�$�ο��$���}�;ʑ��+H!�3!��_��+R[v2�I"L;v����L�@�`cAyy�a�^$Gb��-_���P�m�~�J+����� ��	��Tש'�����	�M�4��8�4N�:�$�-R<�E:����.�a�>{��2�47��v�X(�i�$�jl#/�m�W��6PO>T"b"t�Ni6��ڲ�����P*rL�2�&��-o��<}�/�������I�_4 �M%b�_ڳw�@�0���O���{O�<�n.f��'>Q~�d�����@~���'���5�2�:��$���,v�~�V��=�t�^z�<��K����/����x5Ŀx�f��~	���[� �N�kN�;Q����~ J�]�*�b>d��5L����PnE|�L��7|���y����ܯr�������8��nB՝*��g8�t�C�i��o}����+���o�x�5.v�_3EĶs¸C%�J��6�u��"�8�m�&��m'��/���ŗJ�K%k��R����Oݟ���k�ݢ��:��r�P�rsO�*���гb	�6��@V4��Z�T�~ƕj[q�l�=={�1�q�����s?�s��ʅ%*�66��v%�?������w�Sw��,x�/�zyd�׾x�s�G�����E�B�vʽJc�܋ �
R)��@Y�I��`�(����CDs�A)�h�R$���S�J��{Y.7h)֌#X��0��@w����O�>U��ɔCls��-�U^��'�;KY��o��|����*C��W�&��%~a+<���r��G�9�����R��z"v��AuWe����~�_?m�V։NcX;>>>Ć���>��%�N����-���pC�/OdWi	e�U&��m+��U�;�5|��� �eC��C����L�S�?��?�����}eY</�ԏ?d��Ε׽�Ay��w���@F_I�JB��g���sϓ�v9{��������;�׽]��{����S�EQb�aѱ�@.���^6�TI��I#�^q�(��:wȼ�L�k����+�n��JK��bXW'}���h��\l������,&ѹ�!A)�OX���:t*�-W�y{��#�!u��Y?�j�4���0R������Ȇc�l䷧�?�����iy�E�ݕo�l<��c���u�eЁ�̓��y*&D!]�+��,T��Y{T����'��`0�At7DR��:n-EN�"�|������h���"��eq���r9ľ���J!z˃e������/3��s��+���2U�T�r����}��W���ʣo{{��O�w��@��R9���1؇c��:݄/�ϲ�zJy���j�7+� 䅀2�X�����<E��k�O ��K$�ѩV�J!P[��r��st��3tVz�Q����tF&� ����w�� ���O>^~�;�o�+�"\��)W���8�?�d	K ��[}9[��R�9� �=��Qu��\$峝�#�A:;"����n;�p�'+ٴ!�hñ����j*�[�Ҡpg��X������ڢDuO�/�����o=��J�2�Y[Z�9񥨹(
,)Pl�F��h���滩௨�* ����Q�����n~u�M��G�/��/���/�}�S���P*�"�3�z,� ����xac����o��R��GˋO}�얃"�#�tVHf�?^o��o��x��c����O~����rm���9�0˰��{._��mNf��/p�:,0��#�N� ���}��G�ܼ����"Ew�ɖx�G�}���(���,^[���'H��R����\9���{����K/���e���f�{;�+�_��vKݸ�\{m��b�{��]}0n��K�hC;�vf�-\4S�D�r�vg`�yWܽk u��%���B6>;�~dİ�Qq�Z�D,t�ӳR��t7^�B)2�/Q�	A25�.�p�=����c*<P���"{*����}��������r���${T��:Q^ϵiKW�_|�\�t��G�Rϗ�\������w�w���l��'>R�O��2l�
TR6�rm_Cj�	�$�f"�`cr��I�`sJ��O��0 @�N��t�CƼa�MU�~��s�Pec���7�8�����<Ĩ��������T.(�c Q^"D�An�����M�m <S"�~�T��l�����ƻ��M3��5l�,�z�%G9���u���SǏ��ulǛ})eٌ'���M�m܇�|
�
d�J����nW	L���~�Q'b"N��m8������>[�����_�诔ӧN����sL�\ق�MA=�{�[�¡ٹ����!x�w�G��Λ���Ēa�:y�{I�p 驏?���>�Py�����(o�?�����3_���PP��T`���i؇MV&���
�<nݘ�S��T��&�<:6³�y/������"��\g�tw���HM�����P� �U�"I��]�  vÒ�M&Z�+���7��s��t��鮞�0���6�s�cƉ�`|l{͎V�s*��r4ٹ�{뵻N��I79V��T�$��9���;
�"���B}�5n���5NB�w�R�!]�D����r�r�k���Ǹ�b���(�Oo��G\�F�D����!��}���������,�²<r��p�T���/�0�-(���j9�}	��9&u�H������3��7<ZN������ϱ�jy�=+W9�ӑAhw.��ߌS�O|���o?�ˁk�ؓƔ!$#��a�U}��xI�����L�(3\J��u_���T�������r�����Q��2�F�щ�� J:���HD(����~4K��ٶ]�nڍc=vS��}�9��:���
G��閺��Έ�%�_���.��2�d�X�~�IFD�~E�3Q+ڧ���fX�0�����=�*�13�#1pUO����z���P�����py��'�����~w�+���,z�y˛8�vo���*�s_*'9ox���T��^{����8�����ww^,�Pko�;5�t�*'�,XO������JN�7X��D��{O��������0�T�-+�$�}y�I �`*�d.:��p�m���e	�"�����˧^:_�g�<�,��ѵu ������|�+��D{����6���7��z�>m�������eZ��eD���s1Gd�c�$}� Tfo�o�LV�P��5
cO�*.%�PVJ�Dm�v�ڣ+e�2nW"�3l~I�[~T�(�tDr�wu�ӽ���Nr��;�>����������Ky���P^a��̜bE_O@��j�Uq��c����ڲt�Ry��,י�=t��6[cϟ/���\y�����پ�P/=���R��4���S\y|����tEE�PLe����HƦa-�^8_ƨ��������#G���'^g�u�P��Ti�����,{ş��/�=�)�!۔�%N�ó���
;;��x`J��H�D)���^�j���2TƲ��m�l�L?۸�f�4g��eq<6(K&q8|� ���Z�/�]�`ȑQ�cD�cI�m��ր�6�֣Q$� H����&�:��u���K��d�!ܤ�]�'�\AK�o����_�I����� Y'@��b-i�����sr�0HW�\)/.�䩻�r���������S/���@��*w�3��W��*���xq��O=E�&Fǡ�R�m7bQ�gΔ/\潝��[�	��@�ˤc�fZ��vO�-��MF�g��������֗`n���QaE�C�GϤ��e�tY�4���(��@�m��6��-!3�n��6�Ե�M���R�IħƗ�O��xE,�\y�[��=����7]�j�dV�,��d)�L� Yqu�Cy����WU��I�w۹Z���_�i�*%0uo��-����7�jG��.��|��ϕ��?Y����P.��ܸj��+� ҆�(�E�A    IDAT���gN��P� F@����l��<_��c2:V��\9��ܸ����7�7YhD7YŜ����s�8��H��YB|2��� ��-f�7�\//r"� ��g9]j_a�:�H�J�ݶ�9P|�R�*,���9l�:�УW`a\Nw/]tw����<��LFzx�B9�v�ֶ�0�}����[���]G�8^��.��h�2o��{2�6m�p'�ԺڝTJ����ws�[Zb��fp�����_2��E�xG� YH�Be%(��-��3n�FI�2
�Y�qK�3�a3�,��v��cY��o��<�������/�{ j|D�Zd&33�/�\�>�p�v���G_W^�_^���ǹB�Jyy��ԋ/�3�ȣ0�;�\ִ�"-"������(��DP��I�D�� �_�I���/�/Ҙȴ�Y$N.��s'�[sey�4�i�ʣ+��H�ZفAp��8�wA����͆w�U�-�.u�(%<��g��C�ݯW�_�E�T5���*;�J"���aX��{�`�����g�M7��g������s�v<+�.%Me8�K��=��3��qy�hYrÒ^1��5��PG������|}�xj���π�����o�x(�]3R�&��k�ȑ/Bi�.���+�)�꯳��g�=4���|\(���BL(.�RzՆ�A�oe��!��^���N�����?˼Ef�'���jlB���N���1*娓/+�Q�jV !P�P� �Qv7-��E�t4�.r�J�vt�p�wR�ak�^!��0��p�k�'=�}#�`#��ٙ�m�����b?����8�ߎʪ �
L����H@=�e�-c�7��K����9��� �=ٖ(?Q�5�ye�����?�+�V��?������/������K������\6���Y��s+�<o}�����,�\�x��]��B؄��2\:����{����8�
]f�HVa�S>_�-�)?����,���m�.���֛[������t����%j؜����*I����aGb ��n�!aM���dK�xm���p�2��8Vw�T^=)y�9�T	�ԥⰛ���������(9X�JOr!�s�4���-�,��_��Jܪ��CU��~�'p�g�8]T�Ja5�+m8K�JQR�ǧzt�g�Q1�8���>�ܽ�o�D��f���L9�BϷ������.���P��Y�d���{v��F8�
l��8M=R&���M��a3L ��%"�w�xY��-�ܩ���9�������{�l�E�~��O�i�]��4�#�cJ���Ò~���A�@��ZVb
BB;�xȦԡ���*{m�9�5Sݴ�@n��e�������}��3����zv�dKL��wQ��w+ ,�)w�}���J���BJ�3�(��
Z�A�[�K��V�\���"@b�F)��m����O�B�\
���}cg
����=Q����o�[�ϭ��Y�[ҼMj�x^�C/��j&��\8R��)�t��N�
�TX��8���D'����8ļJ�����7�ȦsP���ǿDIή8�D<���r)?�c�Z�ۑ��wU���Oص�4�x�*�OexS�El�j�ݎ������ٸl��㹣úmno�o��*�\�)�h7t�=v��䬻�J%5�ns�ͤ������4X6x��E&I��V��oL#fU������4��*n��X^gy|�\A�6��T����_�_����?�}(gO�.�؉�؛��6�U�a�;#u\F�� "a�e��]e�F�:�ԛK-���}�r�ˀ���
K��������� ��\�:�&d�
7g��bn���;�����U��;z��E|���N�
��'�/��4S�|�Jt���闝#�m�h���N���a��/����RӖ1萦:���o�D�8��u������E���YT$Wea�2�V�K����5n���]��7��)U��6J�ku��y�SDl�1{����h���r������nб�UlJ���'ʽG�!?g��[�=�L�;o�\$qQ'������y����4���*�S��Ơ_��_-�!���>����j�0{N�fC�A*�{��U��u4�d���?����RA�A�dī����a��#ᚁ�S��_�/q�vl��]w�2������#\�C�����>�����;�(�cc��½��hA4dO����UI@O
�G�@�:dIa�~-(�w%M%�<�T���wѲ�����&�3d�6�����J��O��[����N�����_����Q��F���q��{g&Ƽo|���?����E�;�I����=�����+>>5����F�o#�dס��^���� ����nܧ�;�_B�?��ߊ��D�t6����X*k��$�҅k E��7��j%�r	��u0/̱�K��Wa^�"&u4���?D$�"�m�"y�v0�TPwyQW�iƓHU���ŭ��zf:*�o#�v�$ ��O�DV�qC` ��!��>�8�5b����6I�һDp+ 5��OVl�������a�צ��n~�L�%E�R�'��&u�Ke>;T�3�Fn㛮�<s��/������gΜ������c������Q�ao���zZH���RVH��Fc������O��'�=���(��zjh�b�5�}'4��v=�~P���K��Mi{T8d���]R5|g	���j��������5t�����@�*���c��+����ddן}#�� )���$��m��k�y������T�'�X��[ [�[�e���i���	�L߼�O�����	��O�LO]������5l׸�3��|��T���g��X�W������?����q�i9z�K{R����'��?�٧�ɞ����ܕ�G�h2^ ���Q�`�Jn��d���kOU���d���!osIus�.�6�܇���/�t3�=u�f�q�!Ѵ�Sֺ8�S��e�LYj��!�^�����&�*���^J�' 2ܠ=��&r& 2^��l����[�5~G��V6���t�e���]}�9�F����'91�UV_�����^�&⎡Z9�2+�.���쮄�e�أ�NӼ���_�AӆKs�*���K�);C�XTw�f|]`+?ߔ1è'�mz��[?�ڷj���������������A�^��_䖣�h�6hn-;��g۹^��1��Oee�Z��O]�6f�S��?���xr�m�pZ5L��R��;K5��f���i��Y}�ػB�*9����e:���	}�$F2�h�և#�L�~
�q���!�1�(��[���J�Q:�UB%��D9d�z��aj}*<�/��u�6��2톷�}�DRY��S�j}2�fU�X�/�M�q�(s��Tc�_�r�az��ɿ?��]~���]���s�9�M�mj�gC�'�M	����v�\+Ry�lӫ����/"E`���ǯ�q�b��[g�~:�Ѽ|2�2Mu&��y�u�W<�s�����mʸ
Q�i	��#�a�t��4ܮp����\��D?�������0���WOs����nβ�u��8qmC�_��nW=a��{��͍�9�jaÞa��	7�(`K����j���E�/r�k�q3��Eh�68L9���값�e�z5!0�7Ӟ�U����O��=�Jaz@H�Å�:��L+�<E��V@s*��{�{=�m^��Zw�&�K������IŅ��]%q|�����=(�E�-R� jm���f>UYa�/w�+˨�#L����s�ѱ5Ww;��ѠYN6�2~��]�4�Ѫ��`ڪ��^�L3�kX�Ϩ(f���x�bBX��|v�Z����ԭ��Y�xQoF\� �ET����Ut�rd%�?+#|����&� W�A�_�N��K7����4��^�2LX���Rtچ���a��u.�T��3~WB�c�l�k��9.I��ӓ醷�,�z�!�,z��a#r��{���i6���0�M�[�6�L�����X���c���6��v��H����8ER_݅�0�5A���i�}�P��-����Tְ�"ւd�H1�ʤ	�@�_3?=ʙq����`�K	s�gx�צ��*өY�*�%�����	kqj��%�8d㛶w�YW��uO����7i��g\���n4�x����7�y�����E��dˊĎ�Z�
�d1��e���F�rZ�N��V){M��n�~������~��!I����	��cG$�m#���,O�j��Զ��^?۳��>t�׺ny��j�������<P��\,�3X�l]Av�o������w�K����x=�U�~Z���O�aURݍ�]��W@��5�z?	hv�[;� 2���0;��������h˓ygw��l�:f���i���?��iԑS�֞�|��nYu����ؼ����9��.�;B�=��{��#w��l��A����W΢ns̤O���l��Ӏϴ� �*@������5L�͘]ڤWӼݿ��2�l���DTA�n�'�i��=���O�~�K&�R_+��ܽ�<*�J���O##_ޡF�%V�L����9a�{F;�����t�������p
��̷�g�M=�(s���i�k�$[�9�-�s���޿�G�zJ��n ��Yz_@G�q}c=��d���D6��}�>���ަ���N{�F�z��0�Gu�#O"~���Ks=����Mo0��t�fo�ʹ��z*�U�ƣQӬ��􅁝�v�~���2��oX|{m�{�G�D��2�o<�-^]D�?�q�2�w�aP�7r3pX�!2��^�
V9фb�%xxL�'��*����t��v6��&P��<X�eG����Ul�x�=��|��(�e�X��W�u���������&Ŏ0w�A�Y��0���D����L���MЮ���X�z�q��Td�)��C�H��E?tpHa�k���Q���
��$��4#��tLCjN�F��p���k�;Ŷ��#��ͱ�q��|H b�k2��_��V��-��6`g�t3\�u����,�q�Ӛ�f����f���^�$�ݦ�n;C�mm��,}�j3�f�����6m�m7;�_�׬'�:_=?�I�����^"r�g�A�iH�UN,�_]j.r��s���Sn6v��ٌ���w�I��j\wY	�Qx��-�tEI�_��T�O� p/섉����l$ː�zi��|L�0.�QO�;�2���
�n�1�{�cJ͇�u�IWU�q�� ;T�	wEf9vh,��Qw����6�y3^��()�n�XuO<ݸX8*��Ȳ���!D��-¸hf�m7�)��q�46�+���*�3�����rM�]T?ջ��(�p�9����@�֩qO�׊1EV$ۚ���n�3���~ o B�8����L��Ӟ��l�	t�U5(Z�����ʙ�fy��2�H���8�ӎ�Z��܆׼��`X�Y6�e�S$g:i�-�-4믞f���a�n��mޙ�e�J���
'D�j������M��9��[�3��K7�	(v ���r�?�S(�h`�a C�.�36��į�SUy5�J#�>u��4c�e�"��VM3�l8��'����Fna����g޵�k:�Qӣ$4��1n6�øď�&���$�
�KMK���*��y�Y.�fU_��Q4Dh�l�q�WF�яol�;]:������xN��6B����V�.�zv��I�)	2Y~��l�?���1Ľ$�1b	�V�|c»1	3���L'���>�e���;��} ��Z�X���\.ͯ<K���Ͼ���,Ö+o���ڇ7�7��F�i��=�5���V�M`�/��W@�n��+�J�0*�UO?�M�C�C��/_�?)�e�Mez7�g�,�nqu���ߦ�_�������uw
�����Ջ=馞��D���,QVt���u0��:��I�gx�2L/==Q�^�U�d���k�s���w��W�^���:@��>��������,�x>�������W��=v-�Ҝ�H$Ю��T��n�})Ag�A�#T�g7 �f��;��Yw�A$FS��=�n�W����4#�.�^"{�4�����K�g��Tփ/�a@�{�O�f���Q��mq'��5t�0ӱQٞ	�-����i�/˄~��U1�tW�I�-���ԍ���gߔ����b��Ec<��}sbj�����0�N-���q(*KwTZ t��W�h�[���Ġ����z��O�q�_?�2�l�A�tϴ�[s��b�����kˮ�/���ɊDZ����]y]hD��mm|Y�ɰ��W�.����5��a�M��+�U���8��Y�{?7�΅�?�Fn6r��l��s��f��=lx��wSY/do� ���e�l� L��f�oU�{��V����8Mok�k�8:'Rg�6O�e~鿗^�!��j��d�uJ
�S{4tJ?
����� Z��1�ƿ��G���\ȴ���0�eu�U��G[~��5�>�[{��8��Un���,����"ޕr�_3�W����'O�����������to�Ѡ�B��=+�]�� �� ��4jO��[�q2��3?�f���洧�q��;����1���#�e���龛��o�i�w��nY�����-w�@���rKLZXePØ��*a�s��3~�.˓q�˯�O'㙗��i����f�ϝ;�̾w�����	��kE��k��
|�!� w0m���+IY��-x*+$���<Zq�3^\���t3ͭj�����3��gg��������j�u��#Ы��8����֫Ъ������QM6Ds�	s���u"� �T�N��{�Y��Ȭ{�k��W�����0�����ޱ.�^��4�|jiq�WW���^����=����>=�������{��Y��da�SY��J�_�מH�9��f�V�٪������3�v��~����2L��|�<&��S�i������-|�g�A=����5*��*�}�$�L�6���Dp�2n�SOx���L;�d:�J�ZV�<���'s��WVxY�(���6�yw�x �n�0�����;l�w��D�2nV����;�H�;������Z��&+Q��i'@Ե[�l����8��k�e��lt�i6|�O�uw�A��6�f�QO�O��=�S*�Ր����+O�k�]�Z���&�֎�g{�j��$�l9U�%^��캙��l\�х�W7\�Q_�H{���	s�Y�����[�M?e��؋�'M�����&��ݕ-�7rS#A6����}��\qW;(�����l�[D��$��,�.z�1,_V8�i�_�|�_���5�[�zz����"z�g�5t?����k�w�oöf�ߦߖ!��:�~��b��2d<�7�[�M{�e8�������l�}�B�ޓN�G)�hutz�����n��ۺ�
�`[=t�3o?��s�7�ή��sQ���~Y!����$�}��[ȶ���Z.g߬�ƞ�[��Q�[,w���}�[��j�v�JiDlU�=�E�گ�T����|}����i��km���-��]�i�!U�n�|!5��ȓ<�$x��"6{7�v��*���?w�S�Q�-B{@AQ�����f�x\b���)�t�7�Flg뎱aʓ���Eks��{K��BZI�Ys[�Y��E��2N��፟ȩ�ٯ��m~�� �a3�ަ�_k�<�]=�����=��� �_�u�uk�3n�հ"o *��H���4U�f�¡��u�Z?���7h�=<����|�e�2��m?�p���f��m���2�]�}#w��:�.��Ӏg.��*���r����0{���/+�{=S\�kz-u��ߡ�ׄ�� �5�ifGJ��?�ճ�GW�S"�OC�~Y]��sF��Ou�;jOe�_��q-C���h^R��"Y�$!�w�jm�ȓcWEǀ���`��0E�!BZTR�FV�<�=ͻ�����~�nʷU�J�ئ#�����Qݻʹ��ܼ����ZX^"Sa0�M�����ّ��M���۝T�I}0��(b6�'Rd��W*Py�;���|�o�t��Ӟ髧�z�k��kn�kӕ@��#ߎ�h�3����=t�&
G���Mwqƻ�Q[����q�K\I?uݼP%��Yx�:̼ⱉ��5�q��-����w�����=�ek�{}��5�E�+�K�LQBB'��T�b��    IDAT��W��)J�t��a��=���6?X	�^>]<ä��&��_��i�#��8�9/�7L�aڸ�1g�g��UڝhQ�0;x��7���a�b��q���e�v��j~�
)�69�ۺf9uKs�5J�u�C���ԭ��7�*5�=�@r_���<Y����� 2��O~�|�����!d�M.����u�;���� AQ;z`e����ʳL.��ig>�i�u�<3�z���n�{�=U��v�6��}?��13�uK�L��$�fy�rf�W����</�n�ӭ+,�=�=�gҬ����n�+��B�@m�V�i�I�7[�\;Zys-�t�FW�3�L�يe��̳"��=mȦ�w�� ��d�=��2�LW�H�yj�<#\�-�,���E�T7b��bχt��#巜���s��o8cd����Ġ�,��R��*#:�mq߉&K�Of�6��^8�~�Qe��}h��ݩ �#_k{�L!��ʔ�)e��ŝ�H�E�M;^G���ޱn�*�h��Ӱ�	��?w����V�G��g�c<���EI\b4:��L�K8R��g��ݥnsParb�[1��Z�������A$��U{ �^��'�5�t�-���8*��LO��m�̣�����3�;�J����S�3H�߽}�3M�����Z�#,���_s�1ӌ<��+P�z�I�H���!<1X��b�~v��|��-ի���9�n��;������1J�����Nv϶�fE+8'�@EW��uo�����=U�����=-wԓ���Y����y�n6��=���[�ߍL4�v�z�g����n�NSߌ�.��&G:�~��~�m:m��%�h���sϸ������[�iʘ����I8݈w�m*����L/�;�u��}gg.&�y�6���[��u��-c�ݔ�6�)d�Փ�nF]e�l�Aզi�L#�����<N{���n��,�ni[�TmY�m�8�e��O=㥮{~�z��7˒a���ކ�p����n���f�Գùx�{�B<�kO�K+�vK�u�7�f�,���
-�@^Y�M��`Da�{3�Gg��ߠ�J��e:��ֆ��9Û^旺n��n�{k6ܗ������gڷw���zp��x�յ@��n���.p6zv+�vsҚDG�b\�F�^ڤ��qSE=;Xf����'��Ӎ���CA��e�fK��KoY������U�������p{�w8��E܆���`��˟�r�z�M�
��n�m�*���	����i����2�Aw�;���պe�>�_L^6�z��i�g��~�M�dz�iΰ�[��F�z.��z��{�sl��(
\�ۋ/"�^�b�G=��G���l�ѣ �C<:*��3|l�,��\�"�*$��z�`�X���7��x�q���5L�֚�8m�m�/�l'6��2=���񮤢�u�ޖ+�Gܻ�؆������-�H�{�5�6ˮ�O�yd��=�Ͱ�u3|ύb�(�̸���'N�oO"\���I\q������:�k8��/���,������
���a'$^Gfa��<Se�'`�-èO�a4���n�t�4RL?�gx�v�F�KUm��&-�[�^�;�i�i��:�W�5�o/m<��0J�D����<������"ͮ���[�#���q�r4�a�<nܨ+��}�˼�y��>=��=<���-�l��. �������1��mʱ��@j�WP���w�~-r�/+��L�Y�4'�ɰ��f�m�~m���p��J{�մ�qSe>��Ꙗ�6�iti��ƕ27YGr�g���tul�O��[����]{}��Բꖓ��]���~v�]?���&i��7y�t��m��w.aڙ���'�3�n�;�����
��#�w�l���g�l	p��J]��zAO��f�� Q��ůV�/U�-�f�VY�T�P�3|����7�N�_�q5g|��9�͸�e�2��K�0�t7M��k�2\�����`m�����o�hnå�n'��kuˬ�1^��a#�9����X>�M��/n���=.6�"�8z(Q"'�۩,��9sWܽk��2׍L��e�d�FdFq��fȹ-[�z���]�X�p�,��Qw�*�����ӿ#i�m���2�id�hT�����|0f�W�Q�Y�^i�ѽ'�Q��t�e�p�QJ?�CM%�u��xY�t�Mw[���W:�|5e��{���OЌ�z��G��=ӳ�!m�k������"t}[�����k�q�[fW�C�܎E>�ޟ��*��Nպ�Ӭ_��ά_����=��O�i�kW�g�p�~�=�w)�H��R��}��F�rd�3��gg���ʶ#���D�����L�g2�G��+4�����0k<���ӽ ���O���D9��rAG�ۓ8�F��~w��M�y�A����K��6��Q��݁�V`d%�0VZ5<��g�3G{-�&u�MՆ�M{���n~�iؓ�*�ɖ3�o���~F�>�^c�{��i��M�L����'z������4Y�V7���Q���42^��h�n�4z�3���Twۢ�����ק�y1-ٓ���a^;H�f����FnX� �vS�h��?�k�kX�Y ��~[)����m��j����id2�`z��N�_v�to�[��t�\9,��_��q�4�U���j�Y��ph�N�֭5g�t2�z�k"��;�x?�3G"^�P�|ϴ񏉦q�s�fN$��m�m쒾��o���2 �L��`S�*�ʡX�D���pP�D{��=�5n��j7��~�3�t�3�tO��z�%�ʔz��x�z/�@����3�i�{��@:�q�+�n��-�3ʹ�H�[�4�f���fôj0\����a��+-a��%�HBҦ=�;�����b�T����\RY7�D��������������uvj�r�����:{Q"wL$1Ǎ��f��J�f�iO�hn��9������z�@&ͦ�*�2^��a�r2�f��z���ץ�i[�Vq��gm�i�����2�F�c��/�Id8�/�Ro��*����ZQ�t�,G�A��a�H�t���(o'H�?�TE���p}M��Uԉ�׷���?�FnVע��1[��f_�D��l%��d�2��,��7��Jd�Z�K���6�u�������܌�j�~9F�� \�z�x���ȇ��꣓����i�X�t�Uδ���a�׏��{2?�T��nm�Z����F��bF<��Ong^'�+oRw����6�ʜ={o���	&FK����Y
V��ʒǧ&gx�Έ���1*a���2`vTwx�A}-���2?�TO��t�J��H��3���;Xh8��f@��Xh�$��<��Ꞅ�x�c����:g�U:[U��^���"m��(ʟ{҇�q�$i�ӮDV��7yP�Gj�sNhp��/ab�=&���IbO�o�n��gE���ߠ��>��-_z Be���򧍓���=�$d(5�H�ig&�˸�Ty9�f����9_QN��k �P��3(�\[Y.ss3e��R��ˋ��G�����́�X.^'��|˷�?�_���
B{�(8>�$�ն������/���g��BL����"��yx@�R�N�\MI��܊"�e�N�^�.�:RĦ�zv$�]런�#��.�U-�zp��R��_;��٪^x5�w����Ӊ0]�v���#�|)r5�l���8}�5\~g"�b����G+
eST�'�VWI�SUJC�p�@
���HD* )�x� ���� vT������c��'�b�d�
o�;J������Җ�$�v��\��y�^N�{��ݟ��r����Ʒ���Z�g���ۙ��賵�X�\}��M��H[�?C������~�7���;��<��3��C���%�����"8��6"Ј��DT@���P��H�b����L��4-B;B�
�Jd.��G���X��[=��ꔐ��#3�4(�%(��a�_J[A\̹�p=FDPj����H���r}/EXB]6��xfud��E�j��G�x�2UT��X�A��7��n6z�3N{�~f����޵1���W�W�B{�ڣN33�m�J98;Wn޸�9U�\^ �7���گ.����<��7��Rϡ½-Q�'?��e� �mh�^�+C������,��
^���[������ce�ȁ�|���?���W�cÕ�1oG�d�qU��傲p������:�fWg�1�޵%�G� }�g��lͫg¹�h�F7L�ӯ��!�~]v�e��#ZO5�^��S���w_�ϫ()9v�X���ꐭ����`�7r��e�Ҏ���C��#��7͂����S@:+�[y�k+�@ɰi���q�EH�D��=M^C-�ٱ7��9�������R�n)0/_�P&aU�a�W�ڟ/G�,���@�Q(�X����z�*� \-˜�C�A���g׸`���h��5̲7 �ƭ����{�3��w������r��8��d�yG�/�o�*e9G@~_;Du ����o��� {e�R�@�h&�����'�G�5���7m�O�F���_m�l�q�)�!��1���F��N��B�l��������\�w'}_����������$������G�`$�L�F�2���-��#���h�
0+�{ �:� �v�!|�����>׹���ި�5�y���s�9��Ux���J�k�W
Ѓ績k�|�w��������׃��v�
H3�q�	�h9r��L"���%�����8_&� 7�Q�����́p�E?u�^�|
~��B���J6�*����4�NԵ�@�pՁs,���z
gU�b���֝�f݅M��]2�����_d�D���i��e��-ä.��ٷ�5���_~�r��щC�N�6+���=:>�q=��9�l��y#ޥ��y��Y���n�VJ-"��2\�����}*�q�*�@�|)�ʗnu�[D�0ye��0It�͛ 0�~�W~e����r�� �+\�?_�^�ä�~yy�LN�����ū���	�ݙ�aX�_�l��
H�y�3X�i؏�7.�q���^)K7��[<lt��da?|����{cR\�+���X),�p����p�}�jV���]������Cs�^=үI�~��ԺB��Ʃ�4�Î�e4�NI8Uۖ�v �;q�D��U�2�i��H�2� �wQ���/���wY��q���o@�W��V-)��[� DB�.�Jo)PV�F��dD�g8�2l�Y"�@k�䷕��_K�"��[����_*����ჇA��r`�`y�����q�M.i��ˡ�sP��6�a�౫:�/߲�K$¼��Z��)K�܌nL0�X}���t��\�l��ó����ꤏ�����e�NW[�"P Q :YH�QN��ȦN�D��	�M�
�|;'U�*탰�=ag��+͉�3R�'�[�^(Kg0_��{��c�VWE�*�
mż|�Z�����ͯ�X�����7֜Q�ܾ�><�-�D �t\j��������k�ʉl�J����D����#eowUk��,���QB�%[Q��>6֟������[ʛ����	w!�'U�2�E���;EF%¾, ��ZE��X�>�V�ɩq�?T���4(�fsk	^���n0�^.�`T���T���(������J�VaM��� G�B���+eb��:���L��ӫ�k�^�� `����#�^�nP�32`�|y����R�P�	�w�{;n�)�1jG�B�)Ͱ��+ݮ�M�]dh�ɱ؆B۫-��rk���~�j���'w���}/�/�]ʷ�l���^�5�j"����* ���q�̊Z)�KU&��>��Ͱ��d�Z��5|� ����N�$�ȑ#�sD	9�,�d,��������<W����,��+י��bbe�7���2A�SIDuK�e>zll�k X����v/��$�-�X:̱=<�F<�G>;�oxd�,�|���C����W*7�/��).��^�%�����Ab�$�� �R�	���K�΅�=��������O�M�����m�,��(}�x	�l?��	�#/�vݢ�;��a"@'����o�Éz� 6�nӔ����	=���Lp}_�}������u�n3���8�r+G����iq��ʷe�0�%b'�w�%�N��_��]�"�i~)��q�A)ȱcG�&qR����K��`�u_����Ώ� �*��X*d�1���< ��fw�1�ff�=�,�CJ7_+�P���_����cz�S%���\ER�� K���,��vbb::���f��*z��Dy��3���.��(߶����Vοr��Xܠ� -�.���9ne�E��x �λBgr@I>��6G)�U�_��#�}5ؑJ�T?�;��4���ILG��໵�YK�	�1T��<R�9Gn���m�.��U>��v���ܣ�ܨ�bi�.-l�,��������e�,`���+ ��'�&�G�L =�t��;�2h����b���PaYCj�p��bʷ}۷����{���O���z�I�*7v�ƅ� �K�  �敠֛KP�eq�2io�C#1Y�	o�L\����,ȸ84�����3����k��.W�!����]"��x��2[<^>���r�)�p�K�{(�ty��O�����Ay�%��	D�W��,Ӂ&�8Kt4���I��� K�D6F�4����p�3L~&(r�%�U6ݴ�T�q���Q�j�I�쬟��B9s�yF�ҥ�V�B�6�%���T�zcD���~7�xR����;����5��m����Hs���ƌx�V��~����0�����wѝ����}wy����C�'�]���ϰ�a�.�27;Ų;T1����-X	d��S��˅K@d�h�B�^,�K���k��LM��	5�Z9vN�'�2Y����30cS���	�1�
�W
���������˗��O-�_\�,o|���#?�����?\~闞$}�X;������M�׿��
�p�e��]�1��ا�����=H��P����v�&��4�t����6��{/��jbb$ؓ�����c�������;��ω�R����5�غo᰿�E��Z�� �պ��
��h��WO������ęu�y�zH8(+���޾���|���E�9� �6����|q�I��R�m&��K��U�����}��O,�l<�LM�Drb	ȑqyB��$4
��Mf���,)S��U`���H9��e�ztd�:2�y�tf���rz{�{˵��'˥k����ϗ�O�����~�)��{ϗ��?_�|��r��[�|>d�#�[g ԃ�bP�@�mR���RdV	����?�t�v��to�N�ȡ'çn���/:�fG`�\�9~��Ёٙ�龗ڽK����"���6��GJ��F�xR-�8+�%
��v�|\_�d�������^�5�F~�b�.J�=��"�
��р��n!~��^`�������o��߈�׮]e�u%�k]A\a�bhg'��B��SS6�|y��ϗ����@��P�u���ˡ[�c�����/�O��2;��n���V��C��3� �#�����K�0l�ְ��B����ÓX��?�X.^�h�F^�j9��d���PN�:Px�x���|-���)��jm��I^o���<�TVJˊ�C.�+��K8���O�JJ�07��F�N��btP�^۴v��sd{ն��:e9��ٮ.�u�p۫�o}+,���q������=]jw��Ŗ�]��9�$�r��=%��\[c���*H� !nx�^�V�Ъ�c{fcO~2��4�:H6��-[��tӬLԕ�{�9�$�����������A�X��K��^�>Ϟ��@�nݼP.n�օ��z�A<�ݤ?��>�b���mxk�q.E�j*C�Bg��iD
���Q�Q��%�5�F�xG�D��sK!�^����F <bL'�k[A��M�-�_x��tu�����v�E��嫿�]�G~������b���v(��P16H$L�������4'��`<����@���v5|�W�$�팧ҽ3�8��O���1��/����O?�4���&DV-.$l�    IDAT7�Qw��Bn��!����6�׷��s{)��8����%� ����Nܤ]#s^I��w� +@ԿҲD��<��I6yE��[dB#*�0������|�W�BT�P��Ef�B^�$�}쭏��}�/S�C��rm�O�[\�R�ͯm\�dM`?��k�W���4���H����Z k��3T�m��^+�ť 9�_�ޡ�%S��L[�md��/ D�Ed���|��	��&c~����jϢ�y�b�
s�f�<�j��_|��9�@y��)/�|�|�w~My����G>�I�����h��r�nHV��I�Wa���"Q$�� �A��h�!��/ʁ���eG��l����0�v�hGe�T5C �-L�9U	L,L5!� ��Y�gy�u�,o`!i�w0�{����)�V)����{����x߀2�Z�Ae�+@�Lu3�a��HѦ��җ���"�R����d	��;����W�ǿ\���7�^���<�����Di��IDv�`]���\������TtrJ�(֣��O��D�I\�2�j)�TR�ӱ���p:�Fa��E� �,;WC�`ǕOg�`�Ō��4�PpxP|@=Ţ��`��W~�V=	>5�uc婧?K�b��C��B����=R~�_�kF�U:�WaGY�B��(����Ŭ�*�M��������n����Źb{�v�i�������ؐ�z�¤Y='���#���xrr����ȹ����l�r�=��мڕ~ƦG��:$g��Z�@�[��_tW�p��pȬ���6�65�(���I>�}�(��Y���������+ސ����(tc�=�P�!�|�������XLaG�6K��K���@Mi�\����mv����bI�JLR4�Qc�� �e��ENp�ӄi��CL0ch��[��~@�qS�����(�<����a�S<��j��	�㾧<��2��������b�|�����n��-,��Ú��P�#���[��&�3$n�iɭ94�խ�TY,���Tݶ�.Zk�^�t	q���[�u�vM�	Oɢ!��ms˦���go�/����B3~J���ۊ�ږr+��u �9U�ڳ����Tm���N 0� �z�F�ڊ���1{�,�C�>���'�xQH͖It��H9�#�^�Zo,/]`���<?0 �+�L#�'�v���7��3�dug���iT�,ӆ�8��Hi��r{�4�> 9�:t��A��!6������ �=Ӭr��3�З����3��3���}��{���CgCl69����+�����}nn��c2d�9��v@$O
CD.1��N�8�Dp�+��K���l�A����3�4�ܵ�\���M�Cح��.j_�m�ԁ&�˭�e�-����.��Bν�[������+�� ��B�X5h�תL'(�'�M�ೕ�L��</��	�x���]����!b�q�z�7aC�K+,��h�[�_)����ي���r-�C(#�U��.���1��T4� �e	��[Az(R�.����\�R]`E�.��4H��q�E7y�j�+��A��l�f;�Y�|�ۊ��cL�op>�$�>T�y�Y��\�?���ןe$�����|�ϰ�q����Cl����Z+���V-azM5ipy�:_�A�{R�����5>�̿l�a�)�S��N�$_dv$"��!N�C�&�Vc�s����c��L�븳���履�[��kkt*�?P�A��Y��l�Y�;�m���G
�)�×�u��={_9{�Y��c���D}���[�!�[������^ ٖ
s�r�� �Jt��a^�`�]�`�%V���n�YCN�T
�������]��9(�Q�8yb�r��lh� ����q���g]�f�<�@��Nv�z�_D�93�\v�i�V�)�jy�u���˧>����������{��]��O�83ð)�#�&:L�6	�
�7H�c1P��S�Vm��aj�D�Ԡ=�S��6V��e9c��+��`rw}_�mRtFI�⿡���IVo�T�� k����*K���	���H��2�n��6%����
�c� ��~�`�{������C_em���|���ɣ����x����]-Ǐ��� �A^�^Y�H�r<�emyj�r_�����&���A�`��g��J#�&��Ll�E�>?|�<�0����l�9��d&a��H+�;��/U��}Q�1)�n����r�=����R�EʽȹN�K�^~�W~�E��r�����g�/�FD�u��1��G
U�O	��	e�~�)�A�У�$���� ~v��U5��K�V;9 [��&�@I`�V�bK6f��N2A�z0��j�����2T�;�(Ȗ��ٹ�J��Wi�a/e�2n@7�v�A�o^{7�n���m��w��]��q���ny��s�M��͛��~]d���ؔ�ؓ�����Ԙ}%"�Ag����xk��D�Q/��	����@��5 - "�<�,!�'�0;O�2�2���Wʺ���A�Aٙ��\��b��F�D�׺���;�?�����'O���y�N�	������g��\���O�/{�1ح�����l������BS�6"J�P�%��0���ٹ�[\/���h�ʥ_�U��/�Q����OGm�%y?�q=���V`wvNLL���
��j?�=�6��6>��uxt�R�b�ZY�1�L�����iΊJ�����_]d ���gxӏs�l��a���a�+��?��7�7�K�.���W��D3l�f+L��6�巼|��K[�� 0+�na-HP�An��A
��v˪�j��ǐT�pCl��)����J�n˜f�7G�9D}-����H��������zZv�1S�*�X�5c.�PQ�/<:ʊ&,#�>�F�*��:
W)'˛�t�|^�{U�?��)���}����);{�)���F��8Ƥ��������d8yn�t�m���*[8&ǘlW)m���VEےL?�>q�6O3�ڎ��z#����ro�d�2!H�7�˽>19�@��[2BK�l �Df+����T@�tϲ�=�t��i� 5�圣���ه�._�o��U'�L8���q�E�tj�ʱ�ocY�ɛ[W9�H'�7P��e��|TJ-eID�M('����[ 7�?1q�L�jx��Q����9���|�uB�Ȧ���4��h'"q�l���G�iE���0�\2��Od�����l���&�+�`���3�:u� ��O���K�g˻������?^>��%��
�?�.���#�u"������L۔Q�"H��"L��8�X�g�<�;d'�h��,!���숬�5��?]�1+���Ʃ�W�F�U�U�c�[_[�➍z�����È���,�3s C��9j���z��k/'�256?��ᡃ�����?��������Œ�R MI���H��1�ZE|6��P�FL��s����2�]O�ț���~%�0%��h :.,�v�!�&�P�9���a�Ρ����|�o\"�u�27�-r��$�I��ᝡہ\�h�\	�"� 4�p�rJ夤"�R!E��`;:���Y����p�C�3�����#�R������Hy��G����-��g˯���('��|� �#�#�l�+�9w�lO���C��\�T���Iwu�@"������ҏ��Re���4�𖧆�hB��Ǧ�/��?���e��*e�d�}��%Ûc�l]\ZdQgh��tH-X4J�:[ɬx">5��GEDvT�	�~�|4�p�p� �,�z�;��w�}����G�S,\�����?8;�􁳍����!6(�k�8R�^������HVDn��lَ*�ˋo������,[��{7�/�l~��+PQO�ߢqq�L�4��9 �@9��v)�&���v�<e	lt	��nd�"�Hb'=��D�ƗU[^�IǞ���eo���R9{��r���m_>\>����t\&ǫ�����_G:$$�rұ,�Lě��S"o����v�uwس9EX)w}"����ϭ���2�(��Gۻiz\�y��7��^f�X\��� o ʑLɟT�r�����Rɯ�H*U�X��J$�J%)W�"�P�%�e�%SV��bDi;I(�@"@ �%,vg/��s��f�<���}=�~3+���y�~߾��ӧO�>�M��^/�v�l�;����N�ug�;.�C�=�<rnfn
V���2�`>,+oq|���o�S��is Lt ����fD��}za!V�V�n6O�	��Y����[�h#�&�y�[�]��<�6C�G) P��w�GG<�*2�=��x���恊Р�O�@�r"�}LdQQu���@(�@�J����[h 2A�Go��6(T$�8Ÿ��9׮�-��!��<��F֜��*r���Pa��%��ҽ2tO�t�?`	R���5(<�O�m��������	;�|��OQ�s��=Ӽ���L!�调�0l�_;�4�N�{9eU6�N�&�r��A�Ei�il۳t����=	�,�����ᅭ��y�fL*��g�[7�&�ve(�>r7�m����oݞ��_�=y��=o@�1H9kﻣ"�X{ؓZ���Q��}2�^��ȓ��F�?��⥋ͯ����7�-���D�}%�����NN�Dd�-a��6,ɶ,|�{Qw=�z(�,�|-lX���EU($ϼ���-��[��a�#���\4�����8���
����.�Pw��N�ha��Q��6�ґ}:��OE��҈�R��J�Ο?����u&��P�]nn߼QXf�r�?����^C��B��<�#TN$�X��uځl�X��Du�~�v~k#�滶�8n�H�L'ڟ�E�dh�IVlmK;��R�c3�<G�c!�����ѱ���	xl7q�"(�h�v
$���D�9���`�2L0� N�6�x6�1����ͩ3�l���|�cO7�}�2�bV�6���{�E}�j��M(8�W��(��E�Z^{���Ԏ��!���@�eA��	�ڃ@�!\�)�r9�t�?'�P�-v��A��;�Zw�GAN�[	�7uDh*��@��HKG�C�$�K�и���<���vXҢ�v�P�%ٛ1�?yd�fd١,7o�`)�BP�˗?м��nsE�S�G�� ]�����Oތ �UF���Wʺb���SW�;���*oψU�r��,:(u��P�@X����~�X���";la(��#ͱ�����橱����m<������v-"V�X�w�8)p �J� �t	�� �~��,t�8����왳h�-�󆼝�a�r�Qf�U�����/��x��2������Y\hΜ>	�w�!_k�o.d�SdJ��)�cL��/�%#��l��~���8�A)��.��qO�����K�]�Q��r�4)
�v4��è�dމ�������K�c�騒���,�ad��],�.4o��Լ��+4��|ꙟ@\�d����`�9�C�k�N��v�T�إp��X?M�����^��s{�eJ��[8��H\�3���<Ta��{RW����0�Bp�]Wwzjj�=��r{�ܹS�� r�bpϸ.�R8�,���r�n��}מ��]�H��t[ʪ�H-��N[����� �V!�qa+XB���H��,γ�`��.��;�B	I^]Ʉ�>�urj�F8�t6�~��`�%��f����; �c��P�R'T\���F79�O��&�j ���K��t��u�CV����+O����� �n�����:���������&@��S�2k��.�9����=�D��}��?��\�4È�X��g�h���w`=v��'O7�,,�09��pb@�\��{ �m�[>M�A!FR|�=Qd(�3�H�J����㢻�p�3&���i(�v�8u�D�ХL�K���s+.X�#��� � s,�F]��eK0F8Df����3g�R��8[�اPD7VD���"V,�
�����6�t�h���z ���~�s���.E e�#�@�[��i"� *�Y �P%�(ťLPKQF���(ϩtF^��E���s�߆�B��6*S��vq�C)Ï��l�*utW��9�;�T� :�?� ���v"(7��23
8y �B4��x�?i���n��eP"۲ƙ*� ?����ls�6#�D��gcʹU
1���5�T����=��o�y�Hem���2;'��3�5Ri;��̢���s���T��⋝Ev��#��t�g��Q5:Jav�)>α��H2�,#��q!5�EX+��n.jԀ���E�|7��J��|+�8щa�s��_�p���[��� ����w�fc�V�`I�*�i����9���4>��{�ܹ�w��|b|�Oā�kk���e�1#���AY)����Dh��"�R�Clޣ��bv��<�vG�<�n�ߋ�Zg���OJ	B0B!���F�d��S$'t
�-�-/��Ɏx�2�_��:2�A��ANB-���6�Bn�����D\��2�n����.�?��E�9@l�[7��G��$x��ӟ�bt����DsJ�����@@�h�� âǖM�D�a�>(C�=R�3bL�����6 �N� ��&=M�~7��{��C�C�2^�� ���ab��U��,�#�6�?3�s׍TT���A�">*�p	�G������˾� *,M1�3��B�-�JKm�jzuR�P)4y���a�SyT����OY��Ő&~�0mt�B-V+	�>��&:s�@�6v�F[��03�����2Ɗ�"G1{.�;�pz���a����˨K;ʘ�dގn����h�Kw�i���u1}�vd�7p�#v@�}�+I�m�ӧXu�И�ixD6��:�.t�+]��Q<"���6(n�"������X +��P��6��ɰ��nCGÙfĜA}�s��|��*��y;,r�*ɀ=��4�i��md��6�G��eؖ�s�
�����	��ὧ�NCV�:�/*$M�3]<�`X�`�����*�pQ,[��ٜ�Dը�ҋ����T�z�伌1Z���Pa�O�Ex~�:A˦�iB��N�B���O]H����	��zz�6_�o8�������Ia���Ňn�����z�6eW��ZPT�m�)
ʻe��R$�)a�5~lߚI�m8�}l/������(Εr{�T��4��A=����@ü���,3�2�x������z�-U#�h�~����)ݲ���t3��O���5?��?��;ɋ�L��Q{��Zmבּw=&R�`qup�����BcE�@n5����O���a9"ɶTY��O~ԣ��aQT��p����ގIY��A	��^� �E|'� �!���E�^PVQ>\ � �[�-�CG�I)��0��>�(JWv\�"�^;�����7�L�u�F|��ð%�1t;�&a#,��'
T�DhB�����[�M\H�D|�h��=�Ay�˗/3�,2��'�Rn���Ly�١8|,ʽ�>�a�/z.Ƚ��||{k�}���VB"t��pZ�Z�M��=�Ha	��1��=�я6���3���po����!��q�0�Yą[��LaK@n�;(x�0�LT�%���F��&��p���d�jN�jr�4$����u�=�L5���!m��=ؔ�oa�L���f�!l{b�8N�4�$���AVo<i�g*O�\�4"�=Ԓ%7O{����T�=�y��ع8{�Dsay���'�bQ�*�֐�й��`�P-���c.Qnʐ&�F�5�1N�ܸ%���p���Ύ��,��jwr�B�*���kK%#��?�b�����ʕG׸:a�.JJ ��ʘ���!�d}a�7+X��˂g�� �vI��[��E?���Φ��=�� Ԁv�O�=F�@L�V�3��'���|�q�ײ&n����h�}A�2��RM�_(f���ڥN"l��#xr���8%2X�B��g.�qi�z�8*��:���u/�mGa~����>ق��#!'VT��7���    IDAT9x���K������M1�I�-ymD��n�Kh�(5uOc[�ư��2���m� �ߺ�"̌��ȗ�x�)��I�]�4�ys���y_���X���o�fj�H��:�a�S��<U�J��B5��wZ��~�kچ�=�����&z�N�
�����;6J ]�ۨ�2�;�t��L�c��<�F[R
 ]��e2ʉ�q�$C ��;\T�E���M'��|�GD��	�=�b:r�m(,��e]��',
rZou��� I�~G�5��Ae<�O.,�)����Uiy�g�i�M�!���z����x^�t�#���QYF��KY�;eK�l#˒����1�������^�o�gZ޶��Y7ꃈ�+�D��0r_C����'-�3[�Sc-g��mc��V+���~[�4~�O�k..�=�I�0��;4���[���"�ڠLJ2Ȟƴ��\[�6Y�ʨ{Z�}�+�U�rƱg����l��.��ij��p��#�?���~[?��~<��'UV]�j�PR4a��8�#��^`���I+�tT#M[Xy��>R�M����L,�)�?
ז'��:d���:�n���5��ER��M����zDgD&�l��<�k	�����<�<{�9�=3) �#3���,C(�`ȑ��VW�B;�/��O�uO�����/C|� ��p|psn�c���m�ڣ,�xb��r'R��,b��%U��5:�*&��o&�ml���{f*�r�ȼBtt�Q{�eѨ+eS��kaUJ}�uһԡ�V��
��>11�[W�(����&y2�
�7�q�t� xAf�&�]�,��}<�@��}v� f�]:3������Y������v;���y}s�;2]�үg��L�{�m�4ٞ��������P������N
�������H��:���%ix�,GЍ�G��4�Bn�t�愸=A@�Y!&/#]�
�,t��<U]�Ұ}D��LKMy�%D� A�)�`'��"r����P蕣4'gV����PrM�#�m$J&F�S��S,��̜�@˳(d-�S�kL:�,�;��G�2�B�H�%{ߖ��c;|�V�b��u�*�)	釭\^�{S'�Kǌ�pTsN�,�|P7�dY�6ʄR��T�<\CSD�mh�&u���< �|9�`ƝF��sQ�(T��z��z����dq�T��{n�.�D���rQnY.�ua�j���Q��#|-�I<��H!�g�Q�oJ��Wu��"�aE�%\+������sS������N���9�do��̈�R�N����V���!�4�+����)ZS�E��{O�����sT���_RBJP!�g墦C��v�����Ѣ�Q~$�PxE}�ϲ���;�<�Bю+s ���X���u���:$(G �Ҵ�@9�{HQ<L�%��1�D�w���	�|M��`"����@�"�rq^��e"��\���$"7Α���)���Xp�����QӨ�$05�ƚ���1���n%���~�"��iҶ�GX;���+�&��:k��Y?�%8"��*{Gy�6��^h6��]���O?=�ۯ���"�˟c!7WS�[2�}@���B�Jz�����i���-i�pk�@Y�LC�E�mz��9�m�p�#�;��3�2��aC^JN��#P����q�O��T�CJ��#� E�!�pw̔��"|�˚+E���Do󑅂eb�9MS��Š���14+�Sƾɉ��}�Z���a�-,*�R4�I~����P�KU�ԓQ�i��M8����|�Evق�U�H!���u5Cm����u+�y�W��(VJ?렟�6C�u7_�P�S`/2�	,��p�V�&*����oR����c!��佽3#s���Cd�H=)�����J�
�h�\|S��~�dX�h���ïMC�ՑHJ�[��I�����I!������*D�[�5�Q�g���[���>X��j:Ƭx���N�R��AS��o�u�����<�X�$�
,��P[Xm��.ۤ�C���=�x��
e�y���oE��Q*4+��z�����d�E(�4��U���İ�;I�����5$����k���MA�lӴ-�5��&�ֈ�Y6���
R��Z��6�z��s��!�
�;���f�>�÷�s,���Do�L)��܍��؈�3�JX1��0"��T*Qz�ˊf"�?M���$҄�m'b�p .�M&9�� P:w���X�	���
��~��D9�wNs�5Rs1�o���A�b�#�Px��{�_�?�%�6�L=��0ދfb���@H �H(�k<��� �;�И�2�r˺�aw�G�A�=�mD����g�=T�\��6�E.=���9�����l��fd픰d{i�)e��,�Ɖ�m/K"�Ѷ�0�/�/�Rw�g�0v<Ag��T�Q��{,�f�&fBU�C�������
[	�O��)�e�Yx���T�r�Y�"��fG |l�U�IF<�W�Q�/�����n��%��G�����>�;\h6o��ȵ�k�p�8�r������ԍ(��.T���^���ə�� ��l�l�=���-T_�,�tz��-=��хf����oI0�Y��E�ogvW;��ߜ�*�����68b:�s��&�ٯ�$���ɤR�Pz�Z�B�K�R��%�b"W�sK���l����7�.=r�(���"G����'Ȳ��v�A'���qwCQp� �Ny
���*�j�0�M�$<i�e�
���ò��o\%:��fݼpu};���3l=��'&f����[PL7��ds�C�~m�ե'��%�E��D��͆�,��] "P�l�b���qb����!l=	m�DD�:y�q6N�h�}�D�g�! ��t$@��b�v����<���GSD�w�#E٥��;�_�Z�؞L$��Id"�cg.X�1�(iy��:Y�tYv�DjY3B��<��wZ��'({8!3�[��H"��д���I'�(ID"�".�M���Em6�N�C�L��<M�a��,]y�E���tg����y}��Lr���&���E�BCxΨ}��X�mt��1i� Z\�����t�̙�K;��
P���2i�Dj�}Ԃ��	���`�]z�] �%��J��;1�q2�xC'�HFܛ(�(��e�<�[�3��w�|�!~�C�~:����O>�6��)��:�����!F�¦�.�
���"uA�9ڕ���Pg&�¬lE#qD��ә��\qRr��M�6����n-sG�s���s�����!?�B'$��0ѹ��"�,�ڞ�!��w��v���Q]	�#k��p-���k�k�vT;��Ȭ��[>��A4��{nl����׮\9�KA)5�B��ݭB"H�L	�����*�NlV��J�F�C���\R�(	?�����6���'��&�����
��^��<����g���yW�|��)��b��=�.�Ih3�����'mHW#�����b���3��ӡF<�RD��66�&(��'�D"~����וp�1���_9�av�֊F%M����G:R��d7�,����D#�(����i�u#%+JF�7g���tf��r�����Й���Ǣɏ޾��j�><�����b?�bY!�
g˒K�h+l�Dl��aie��ݶ��/r�#�������Q���eHdag���\��^j�OI���$�)YT �'��0�FK0�N!��"k~'⚉q}�$B���;�H/��˯��j�/|!�^�f2�Ss��z""�G�y��8�Ȩ�7���킐� �M�]���?�J��m�8��|�=�l^ �=p��86�Q�] +{IP9;��@O�-���䫿���HPxu��=PQ;��шJ.����5���t|�BD���tӌ̬c���G�	������$+bF�Ng++�a�pB�-[����ͼl�|t��iDn�4��[��,v.���(�q� �u�uaA��Cͱ(���l��V�B��,X*�y������N����H~[�D�H��"�)v���{F��k�Qh�YF9��s�8qT"�D��=���8S���)�G-Ȣ8y��/�{��.G>lnrq*[���\�.��c��J��a�INS�2q��TaH��,)�E=[���i@�bS^Ev¬P5�o%�iڐ"�1�4X�@���Q��d��zj�x���v:�2�Sd��F�&{�|9����qD�)�Sq XM9J�E2�v��ߦ+����iٹ,����� X�#�1�i�蚨#�n���`A�O�ώ}�k_�~����/�؈��9r �m34	4y��:����з-���!�F��H�F	�,���G?�߇Ø�@��.qè�\E��F��C�ú�����`�;��!;���skو�H���TEv����Z�6�o"i���5q��Uz{49�-.�4�(Ԛ�hv.Y�,AnǆB�ccBԫ��2��ǑN�y�ƵAE&^�.}���3��7�BI�O��Է���l�-f�4x�|.�p9ϑkȾ�޽��H��=:����w)��U�����m]�*�����m��A�����L��W4�Z�G��\{����k��&p�
16���3&�pO�~�������HN�ʕ��m�qXȾ_3V̂�XH��́��Ʊ!��&l_�#ņ���$C�p��B)ʕ}n�U��1N$���{��o����b����@!�^��}����1kc�l5c�,{�ANr��JL���z�c�b��%j�/4�����f8Ԓ2�J������FƳj�B�H�Y��]��$L���1��s����G�>K�
���z*��鹛H���<W}�ki�4W N�u�� }��Oe���HZ:UA#�t��<􏼈��mj�ac�t�.�~�&�J��8��QAB6�t��X�vwƾ��o_{��gK�tJ��=��	%����H�I�("ҩv6@ܸ6��2��*�"�5e�K�eŭP��$$Pt�I`�@Я �,�Hnh��v2�ϩ�7v�8ӈ��I�&�^i_�-,�,���'�4 �8ԛ=+���Nܰ���}+w�B�9��MlZ�ĭ
�̞k��c�">���1Z��f��Q�3:��1�$���]�h�.�s	_v�f���A���������߈''�&ᒰLb��l,#*��!,HR�Clr��:��:�
�r*�$lBBc�$[MR����]:�~u��w"r��m��d��w�X��zd݈�P�r� ��i^|����e"�},����l�&�J;�e�c52(ew�I���(��C��^j%�����wm+h:�.)+/�O�>��������i�uD�8c�qG�2�i��V9Ijǭe�"�T�]7Й�à�H��~�2W�^�֫�+n���[͐Rx{Y�l 'i8�m��'E�Y�a2��\���r�dNM{(=��)W������hٰeg��ԒNva�@#�[tB�E"M�D��C���Dh�3��hvd�<�b�;�]���]���e�ܾ�1�ʴ�Q) �?��K��!J���Y�L!����>�^MЖ�E�1M��%cD�n~H"%��K;4ǃ��]�EE�ߣ�Bo������=tg���St;�	�O��a&�J)I�`��/�3L �t��MW��'N�!��NL�q���DC�����p<YR��R�O�3�<y�@WDA\O�b��YĹ��A�Y��G��0�EZn\%z���	��q݌}���nP&�n��$'���<.��&ؘ֗���7���"���z�O���D|��'q�c8�-���xxO�݄(-��L��/\x�y��M�\o�{�&j�����{�`�m��n��m��eЮ��}X��K;�(�En����A����#w��<eD�Y� �������;*���4ul,��;�X�A�K��0�Ҕ�.}QwG��eNw� ;�=۳-�ω�îq��.���#����e{�r�� ��噳*�
���']&�JI�һh�)�i�YF���f%����t��L4; ��Z�8Go��������'�Cq���5;�z�7n�'�ބ䅎�un�ȭi��'l,O"xڲ5�s��"����4�#��D��
���0v��\��{7��Kw���*,���e�q�0���'�k��Þ ��&�L�RG����x�u�4Taʸ��-��>��yj0����ԩ� Pgd�ۍ�!�7�m(vQe'�T������~�#X�'�7���=�
q�e�k�{����/��x��AMX:?Ź�#�Om;�����C���A�\͖b�@�ゎ�x��=�_��1��v� Gc�$��l<�i~���܅'(�"��,��:/����K���-�t�����x��=q���S&�Ym�ʼ�Z٨B�^�����%�;B*ϟ[�0L�)�I8G	�Du�٠�S�����^��d,�V�zu;�%����01��k2ϴñuO�l����گ����:F����D���Q��L䎚u�RJ{�l	KڻF�
%:&E ��<�vR{�`��J�{�\)�yd��|� )��a=I��ׯ4��+���]?^��ȎA@�)�HƩ���)��EV�r�U�ˣ�CΞI/��\"�N����&��ҁ&Q�:s�C�Ň���с�&�=��N$�l�)vQ���E��J^�'4�lA4OA�A��)7T^�[&a��	�ω�:��c���(��-�ě�B��,�E���\��u�'$�� [�������g^i�-퀗0�ɶO��6n��t�}d7�ac1�bw��q�;x3�I6��8�b����]A�qVJ[	J
�u��v�����k���PC�-��I� ���Y�ҟ�<�@B�1����R����Ypmݥ{;�35<�7���!������-4.
���3�ܭh�[(qp�����in�@j����̙����G`�. w_�p� +�Fބ�g���2���(����I�`��A���T<�]Qc�t��X:�pK�y��bP����^$B�c�v	�����F��]n_���_��n��}��y x�N"�j�R�x"��O�_�e�=Cg��f'K������c����ܑ~\�&m-E����s����-�$)G�:(�JRq�e��J���iO��)Tի �ƛGX����w�0�,�m��Lە��).P]8��p]V�:�x�'TV]HPT�[9��m�R�2V�����P�Y�!��ԥ��(
�&O%"'O�cO�9�=�*��8cP�R�LP�<e=�-�,��D����}�(,���r����tA*�^Rm�6�x�RH��޽׼��͝H
�w�n܄y�$�>�A��m�aO��a����������.>h8oA����?_�#\��I�~��]�)	��v}ksdyee������Teu�P�(��K��Ah�}46RK7ߣ��y(d��� �&���8�`���mv�Lr6����_������]n��l<��T�q���͛���d�`d�f������tX�������[Pl:��_"o��ӳ=F)eA%�;exa^����Ű��&�1�.TX�ؠ~ݓ�#�|�قUP<)E|��b5��"6��c���;�����)�}K^�f�{t:�J�I"�]��L����Q^/�݁wF¨֓�B3Ǆw�^�YB�}u��3�'������j����f��]ξ��|ؤ�uGsWR!q���V	ҳc���ĄR���m#;�����M*�-��ǚ ���$qº�
�F��]gpn��؍C;GtR�2v�*m<��s�G!x!��,?ίk�jlI%��HNv��;\��Br!�<c�t"�
8���������,�GOn���#Peq\�`$�b�,�믿qՋ�ۋWmt����F�q"�`�2Q,�KB%�xS��MeH�]��>��ʈd�m��2߀L��	��z$�g���P��`Kȇş�i���k6�>�0U4*/^z����ԅ���$���M�Oa�#�nN�U�U��řy&���o4�\����*��YD�w�%Qua����#pP�L��[�m�O�Y�����Ѳ�h�]��Y��!���A�p����KKG����{S����B`��    IDAT�$�KGd������� iGl)|] ��c�
H	|��ss�{ڋ�/��x�D�_��_������.*�d�J!�E��. M@��¨�Ã3Jhԩ�(O�4j�ʜE�I�SF(ҁ�y$6�u��MeP]W,��u�c���;�*��T�{.�w��~�]VI�2�\�'�������c���/a�щ�HB�o��Ǚ#x?���o0Y���5&�WB�	�\���U���f�%�+�/�=w�0�6?z�Zȷ)�2xt�3�z8�Ԙ�ؖYN�k�ᵋt���i�����^U���K��X��mf a���~�ڸ�u\�4``�B,���j�-D|s薌p�[��X�/�`V�(c%2�av_ �G���=V�8�5FDzN�T�w'��?�����w�kv�{f�;�����j�y�y���p>���#���Aᧃ���X.��eTD��E��9�:�DӲ�	G*R���L�Ι�͛Lޖ�X���\� �,�;y����-���D�&�gf��F�;��Ǝ ��oG����`�� ��Ӽ�Y�?9E����l��A�䓟D���%�_e��F���7�T-�Ă"�\X ��>�}
���6�#�!a��#�B�4�s|GmۮB�0"�D'��0Ϸ	G��~��ܴ��5q�QU�h���&}�4+P�6~��)�Kl���cnӊk�SJ3�>G�B��<��1�a;\�@)^��������ɕ�g�]'��<���U�Qv���>Ԝ9��L�\���\�/�
��O���ocJ��NT�2Q%Uu=�oģ��0�.���B�sP�׹���������O��^��\찂��ajj͌N�����4~�<H�d=�s�	�g��v��T�مMR�Gge�͛��ߺ�d���4�$��J���?h��G�1��8���9��e!�Z+C�*mi����|k�//m�t+��7R$�q��?������o�.8�/e�VHv��cϑ���D�,[jB���c\���%B��d���x27�k�f��@.K��жW;�y-������i~��~�;�_�F2.����c�8>OX����_Dķ@����uU��+W���pr�@�=2!&x ��M&a�DXEaqc����[R7=���
��[�IK�7��P��]��Fѻ0wU�E�>�"�P"���Lx������7����Idf�`�k��me���{���Ds��Ǜ��1���kq�<�� )a��JJ
Ֆ ��ؔ��K9�� ۰V)��>Q��i��5�6팧mZOM9�)�	G�|��#����[b�Ka��Β;$�q��s�@��_p�B� ��{g��mT��M��{~g��qU�+����"������ٵ楗^j~�7�9w�Ls�!.��e���1nM�������;�_�P=�F�RZ�xd5,�`Аi%�H(4[n%��Mfb�t�^w�Fy���<+�"G٦������~��A�
�)��Ov��ń�Clʎ�e�*�y�8j�ۨ��F��L����N��Lrw�?���/�Q�v� R-?��&\:�.+��>~�[�fQ���&�}�_�m���o�u"�A܌8�q���ֱ<�!���:�z��݃	�fe���P��]3��&'���4�;��Z%�.�l�"6L�@+���wT���A4������L/Ø��%j�EKJ�a<"�IPT`��r�+��߇R�5���_r�I��	��h�$o�����3)c���U�&���1�EU`OHoTv$VT��fcɗ`h�c]���t6�Nq?��m�+�"����l�F�P�����@4	��&�O��&��0y82��8����VHE��/�ʪ"�JY;,
ua�6`Un����\���B�����b����pM�� ��
O��]��=<�����Pږ����f9��y��h�{~k�)^:E�I��c���	�԰@��v�:7n���d�A�H���~���&=I�����8�>����]l[�p߭�ᇉ��O�$����ߙ�n~g�	�T��!����`=���{B�f�/}�K͟�髰j��j�)U��b2'g��E�O@��X��V=��F�BƮ��j��	\?�LZ	MR�,\��Rz�AK�aQ�U�M��<5	����`���e���K����U�"<)���"���Jʍ���F�A��ڈ.
��	b7��[P�;ȹ��X��<�ؓ�����n�дܼ����F�
�Zmm��� �D���529G���}�d��G����i��G�u�oG ����D�b�fg�����d���@�d��1K�9&r� ������������.�.��̹��FE�� ���țk+淶F7�A3y4|hڠjT�4LY5���7�˿��(W�����g���t����ʟ� +�� �L�<|Q5^���_݈[��;HdV��
H���-/��Eˤa)�TG��Ƒ��|�In9������l���7b:��Ѫ�IY5���z8�U�ue�mpP���EF��\~�-p�nq
6�c�g����;��c�V�3�����_�~����(Hm4H);��'�ز¹�D��k�wS�]A�ҾuZ�ƒߓ�����]��ī �`�u�ub���JKd��=�2��p����u���\�cs�R�_k(P +׆����{��V�F���� 09�G��t�xh���e؈����q����o~���_�c�qq���A�6�5��Ų��<H�0�OOAڛ�ڍ��[�����#x|�e��j<�R��Ҁ��ičmf��`a|��C7�}�^C���
�È`���;2�k]5U�:g��|5�{}{y�O-��1a܃�n�������赟z�y��w`5�X}
9�è�.ѡO4_��>�#'P�� P��p/D����6(���G�z�"ڔ6���9e9��}W�Y����9=kosks���}�2��㗸$`�8�%P��ytss�� bS�ZꣿҔ셆kcE�����n	\��~~��"���X���{U��p����}���_�|�7���)9YXx�	ʇi|ON�>�ô
O(I��w�����a��My|���nj�Έ&6#L�%-� ��XDY��I��$��۰8�;e6�RﭱU�<�sU��]V��p��?�����)�ҟ��K �n���W�h���(�#
꽷;�|��Vs�:;�鬷����0�H-�(C�L$��a$�~;���Zu�8ܯ���>����u��w���V�?k94��\�u�Wp�a� �$��Z�aw������@�IdvWNj6�2��q����E�'��}�0x���e��;� $V�l*]�����H�����?��PM� ��qg��d�ć~��~���!R��<q�,�������н�v�[��"��ܥs���{��Ï����u2����*���65.�c0+G#���]v��`������b��#�A�)ܗ��������1���*���͇/?�&���{|@�6�������_i�M<dg��*K�^E��k ��bC�������_T�H?���@��S3��`���#{��b�)��bn���'�ߎ6�B��N��}�

�Td�dr����Ϊ�bA���N�$�fq��>��ne�����]��w;�(opЄ�8��dr't+
ߏj*���_dQ�f�}_��N����� ?��U��\���w�� ��`'�x�ѧX�9�,]{�Y�}��F��&���ȱQq���1�Un����ܜ��q8.u�S�.L6Y�f�m�5T����w���Q��gP�E�wuce��>���s�.�����h�\};��MM�h�z��t�x�u.oz����E���-$��� f�	�	F4��XŶRN���BJrGP��:�ui;B�ǲ�}K�O�-�<��p�� �%r,�fUdg��%E�� ��K��Or�Eg��lЁ_ܱ���4$�b�'����ɳ�8����������'������PA5�6]P�<�-W�e�(�տ�����w����/5�=�0���i�ns
����mx��P4z�����x�y��[L��u^e,tY������1�%^+�=�W�7�X��;l:VG%�Oa�I�=v����0����܅�,6�o�.6�Hw��B�ݵ��ņ�吜\x��'>
�\�	�[o��|��y��7U�3��H3Ok�+�!�Y��	:�@��p/~���1�*��'%��g4u���Qzc��%�(�lR\�
p?��?�^"9���J&��9r��{���(�OT�V�����h�5\�؉��/G!i\������X���=��6-����d'�A�<� g�"�mo߅M��6_��d��s��<G|��;�������g�����#X�h�����Ϟ�r�zIg���de�ns�]�O��7@�7��;�P��d�9F�	*T� ��1�i�w]�$�ͥ�97C�a�f�+9w��w�xͷ�����?D�{͕7ߎ=�&��kO>�qTw/4/��F�ЅǛW�����I��+�Ҳ�~�|=<�r}�Q��)��`K9��#_~�ؾd;�T]�#L��]ڿ�uf����4�`��fgΞ�=����.g?MЦ�|�9r?�4�>{ʔ�r���w��M-.���5d60̹��@H%X���-�9!Y!�!�����l�@
�O +M�H�d&Y2�/��oTH�Ѹ^�� Sf
+wʩuwO�;��c�������=�9X���z���Dl������c�lC�<�j��z�I����:�\8�p����W�ջh"��iF��<��{������wY�tTpb�̺�=Z�/�5��l�~�4�ف�G{ԳXPt��t0WYY���=���.����WG�kWO5������o�f����,�~�
�o(���@�. ���77?�Uý $��^�a�?$D �b�D��D�tp�hwޝ_y
�ߎl\&�d>�5�c�j�g� I $�ۨ&�)b����7����{I)M��x��V����\����&:�s{4Ю<�%���m��V&�0i ~�ʂǕ����6�t�_�q3��ɰ���>�	.rV��?��4�=�W���K��|��A�����2=�Hl�Z9�\{�G4�Xs��
�p$,�<���m؞E�X[]n�.�
x���N�+�q沼ƍ��|���7���4gΝG���h+�6�Ї�����eGJan/�B � �S�6��� �������lmQP'���f��׿l���s�E.���ĳ��pI�.�sT��m�|�8	�L?ä{Q�*�St\m��nJ���J�s'WkQ?�L�������W���.�n2ď/p@z��)SS,:LN��ϡ9%O�C���M"}��]V�B�ܥ�S�a|���3\�kk2��U~=fN�Ņ�(E����}&�������泟�����[�6���	��� B�Bvj�Cl1Xm3�{�Ή�g��<DgagM{k��?�ݥ�VA�E�G=�������-������2�b�����?K�@T��ۻ�2R������M�o�m�z���^|�N�$|g1-/�Lpq��$��� ܄}��>��/M�g{����SX�fy�V�r����������j;S�̇��Cn�m��$���ڙRc�Q�;3;��qoy�mH{���P�"J��-;���
kk�})nx�?�!0�5	�3�y�{��N3Ͻ�o����ΩT�|���_��|��h��ȇ����O7���������Os��$�>�\��@Yذ�����^J���i�Y�c�P>�L�yy�F�V��MOrM�z�4����+�4��WP-8*V�����I�H��~��0��0�$��M�����	�LL��L� M���s��?�J#,}�,�g�����v��~�6�)�Q��q�¶�2�r�5��M a",AP`�9.rCb�ҫ�ؘ�;�x�^�Ն��1�Z8{f������f�+����6�D쌛��1�_�|�P�W�JI�ƺ��L��.�a�������4���������qs�҅��?�)K���9��N�U$rh�`�ץܻw
����4y��[ל�r�H��]N�e�:��Y��v�F �H�2���N�
+��v��Ύ�A�]8h����2�:�5+�N>��]�Mt��k F
>��m�ap,��F�!�2-C�6)�QM?�p!}�e��H���i	=d�ҥG��}�QD���흲s�M{�ul�_o�_191��<���� A����̘4� >��w��l��-v������2\>�'���M㷏��^�2Uܨ��h�IIfX�t���o~�y���a�d������ͧ?����s��󋁬��PTTHY�]�\ZZC6~�d%�R_ܫ��6��}�.�Ŏ�]&M��W~�n�[��`����}c�C�ud�xY4 Pz(7T�r�	�&e>1w��X��Rt�K�K��#2	����^?��>*�:~�6�)Į�E�I�f<���x�s�ɺ��31={��D���<G�92�������U�d�����I��S)T#T@�Cӈ<��A�d�ׯ��V���'3��+�wӁ+�)�&g�y
�j:�lp2�z(�Ȯ��4����Ss��cPՉ���χ}
��S��4��	w�Oq}��a
EG�>ù��(Tv����x�����U��'Sy��w86&W�pQf�� /�Q9�.&Ċ��g��U�wx�������J���~�[ï~؄e�ǧN+"�?鞶Ά�W/ܤ���izq��Wp��yn9U��ܹ�9������b*�S���A��>��>׹�q �4���B9,��M
��OX)ˎ�
��+j��7�_׿Fd�u��w;���w��v���w)�[X�B��( -+�S�ҽ���
��ߏt_��o5��՟�H���w�g>��泟�,�"�:�3���Yi���&[����f����W��|�w�������C�/����,�c� ����Z�(<=|S�*��Dd7@��(����t� �����O�j��0�:��{�lZ�@{'��.Q9�C;稫��ťK�Z��^\.�R����{���݄���Z��|���)y�0bDj��bں�॒�gE#2?����2X�L?Ӎ��`��1�o��d���H�^P.�
�
�p���&��F�ӥ�<���[���4����������'>��,��YF;�g>�S�3�<K�x�����k_��P޵���p�ɝ8�vV#��V	,�n��K��� G(l!
�,�0RN+�Y.\�D�:֡�]� �m�$���%,¡�1��I?��w��3h1D�tK;��Vit���'�^g0]�HHYB���+W��?����DH���ٳ�2qF�ћ���Qj2G)�{�":�QunX�`"�&��w+#`45b�4��J��0;;�2���"�j��>�hZ+�#Vq�8�q^TF7�za��P���7/8d��׿��X�Yo��E���v���㗛ˏ^n�g	������
[�)P��p��R�3N�P���ɲ���s����������,�c8��E���0�+	ۂ8	'�M�׶���d��=��^{f܄��i"n�Q�)�u$��]�rz�W_�
���G�>Og~d��g�,�}��mB����ۂ!�Ʌ����d�V�D�t��w��&�j���>*|ݡ�8��v�x�m�2��|A��9��*Z�=K���臨5(��G����m�[yEny��^�Ҽ���܉�mΜ?�$U\(�����Y@vl��"g8��e4q� H�+�v݀  CX��C��nvʣL�$��c���w:�a�m�LC7��N�-�
��\�ZI��E��)쫣��L��`#'9�i�d��y�[����#h"���	#8��+�ʊ[�xĖ�|u�֩��;�?,�����LC ��}6҉L�����GbšR�bX���(��qM ��8i�	��Op���8���ltU8c�EG��Nz�	l��RA8+Tٽ�^��DHzY�0�-.u�N:��}3#��*a�߃��}�[�0iZ�������U�C�t��,|8=8��I���7y����
��Xj    IDAT�:.rC��!��C��ua�<.l	��iL�l��.*��U�^p�B�
F�~�>�³�1�^�wV?���~g�Ek%�_�'"_4�X�{���@R'��}��db���pl�"��;&��q�]5"�\��u�#L���HGpC1
X����7.�
��^��Rs����:f�e����0i[�2��%��ݫW	܃��5��6�n�+��V��K�d��θ¦�R��#�mK�A��$�i�C� &L�Z�>#����p ��r���e�_Z��q'���,�O11����դ�~'Y�L�p����a2��K�N�4�b�( :ÔR�/�&�ƙf�a����zxfHH[h/QRB"ew���8X'yIw��c��v �)cn����@L���|!x����zdӱ�=H4"𐟄U��U=KZ������8��{������m0|���OyO�����:��YC�(lXa�ĻKK��X�����m�Y߇�t=hjd�̘?tG��B�;�V�P��+gE|��چդ]��n�դ��2̠����"r�qZ^/´iG�d��3��8�Ӷ���r�w�KU���bCG�n��N��@:Oܘf�uo�.;}�b�JU���z��/U3n*[��-���p%���/���Z�R���r/a�	��Z��l}[�6!�K	�o#��E��N�p�'��K�|L[�W춠VO	�+��w������\Qs�(��.K��ذ!f��V�E�F���%Y|qX��hYP��6�7�a
P�=\��%��|�a2��g:�G����gZ�1J)�u:���"��Y��$k�.�L�,���cޠ��W����S3!
J����%��ɥLN"�
ȷg�n�u��qe�UZ�;ʄ-�ηv�#��"eY�`�i��0�m�.�|��p����o�k�:�~���)�Jx���/$JIHsq���YAv�mcc:�A�G�cSnϻu��������&�����451���'�/*�A(��ul
$0(��PƢ��2'���|�V����@�q(�Mi���+v3��K#c���zR�?��F �Di�2qb,�%,�hU����gWM�K#N���$p����6�Cs��V�o�X�|�쑮a=�d{��c��)BZi����nl�(�W�X�,��9ҳ�i�U1E�,ݵ~a�¡n��>��������x���i��j�Љ�CX;e(�a���w���1=JCMAw>M��nolq��̱��tjԳ�'Bϖc�(����F �S�@2�QS��w��mc x������N�&��wڙ�a��n������_4�bf��W�C؈~OvA�;�+n}� ��2�V�!���8Y ��WsX�[���{�����"��=�h� G~a�d	�`_vİ��3L:SS��A�4�Fn�p��THr"E�%��B`G�̂E#�ȝ2���)��d\W�2��h��
f8��d���4Z��_���S��0�vD�#~I�_;]�y�߃�&�I��q3~���Ҏ|�G�3��3�0{0̃����a��a�s;,��T��)ÉK>���th���0W��\܎�����ds�kJ�1Εsa������-��o�bJ����m��gE#L�,?ϯa���-���`�t7\R��C�7��|��|�ߴ2�v�+ǍΏ�TJ���Y��˸��a���ؑ/�uzu��t"l[��~���y���3���,u��1g9�Hʹ����Zx�)�	b
I<��(g��-�A�5
!{�U:Q����<r,R�g\y0wD{!E��b�nAM�':��}Lô�����dڵ_����+o�1�=���e`/�.�}�_;ޱy�?U��I��G����w'�>��dxG�ވז%��re�>��5�V~k[�(W�Ϡ_�^�G���c�sX��O^�z�K�ޟF=Ac���؅��xo�H��sQn(2eQ���H4���,MaDz*&X8+0ht��{��q�����}0��oÛ���y��i���)��4�3�;�]��Mr3ﶺ�/!�M��@z�Nh�ǰi���m��&���@^��鵟u�poӬ�3f�i�skz���m9ĝR��#d�8�3���IC��d����`��F#	!�\��D4�J$�(o)��}Ƨ6	�t�oä��T��]��p�M��W���ƩM�g����O|ݣ��ѱ*+~�1��">M�a�4�rK��Ԅ݂*.�N��D�M/�p�c��&�yT�{/^ێ��`�m��dX���Bm���������U�:�������R;+m
���0�?j�X!nO��������V4"�c�d�t��:��+ Ȱ.����3=,^ϿM �h�_��[R�K�q2�an��i�e���|������r�wڃ駻v�e�xo�2�`ܬg�>�n\�"L5�.��i)#��/��a��3N@z�96r���Ǣ�x�E6'��<��@�XU��DP����~�DA~;*���L ��v��F�����8�[8���.W��?)��d����[��������=E��k2-��t2l	���ю���6l��μ|7M�i����H�jS���W�k�`;���	C�3����7�u���Pf��u6b��Bܨ�Ɏ$�E�6h0�D`�3zk�Α�ɱ���Z��d�0���^��*JV
ju�����6��ig������8�l��x����ey��'��8�n�緋I�ᣛ͒i��g�h�ϴ�i�y�P�o���"�j;:�v��v�=����["n�Y��2����z�q��u|���[�6�)�	��M00Cb3+���=T'�����N�<�=v�CՏ0�Gnd�/���߂�߇/�&��Ii%!Y�ao��E�(!��[�S ���n���vX��������m�:y�,q�7��Q϶>�!�V��G�L���ȡ�O�ɲ�����g���̑��0!�m=3�LCgœ���x����#���p3n�+�Kăm���%k] �*��x3�^S�u9��t��tmm>�:��C����S�m6Sx+�����(lr�0�%�U�1o�5�"��
����u��/ݵ�=�]���j��{����RQ�u����ښt�w�3���:��w�ӽ�o�����^��'�M/��O�yf�����u�7�|�N�m�i��(�rd�FNU�6�+�=tq��6Ϟ�~�#�q)w+*��A4�%���}��w':N�qA�
ʬLZ1N>�1�,�d��n/�M8��˰=C���U$�&BԈ��ie�3�(i�� O�Lw���5��l1�n#�f�C�^�(s[�3~/,�,�w�[��T�[�"�-�3=��h�w	Q(k�kg���������8��'�i����m�k��N(/~H�U�bB7"�t��7��4���q&�Aa�}�2ԋ#M�GTlaő�n(�P�ر`�Q�'Y���jx�d�0����⦿����rS#���>���du����W��nRk����n��ս~L_�|�4w�=�r�������]{X�_��^�y̝+�Pn��gR�N���v���s�9�s����#��=���e��;r���	���+G~ æ�f ��F����XAW��I��6U�tO��	�L��}ϼ|�͠{��v��3�nX��c��kZ1�gtfq��T����!������,S�����]�A�����el#�n'K��9�N;�{X�u:�_/�/;v6��t�n.E���)��Z�a�����%�%��1)2�dit���g?Op������4CI�m�*�8��^������~[���w�����n��B�=�nz�QS���aܡm|�=m� A�D�*�q#m��zؐ�K~۠��Hl�@��{�a�,�@�(S����t˴�=��'��;ߵ{���Q�v��а<���a<H�F���*�r��ylO��mV�8�]��sw	�}Az8U��fشН>1�.Az?��8;R¤\�F.�4�
r*��JU�|VT$pE�NP�u����>����'�� �1��Nʘ��]SO�q��$�k6@�x��)���5�9=�ʼ���!���E`��{���*�:nl<���ٔ��:.ZT����������Y�D��8�e}�q��x�<��?Îia舔��w�a����$d�ݢ,�u�����7M��<��١i�� N��%:��B���i<`����'h��7�=����Fan�X_��;�#ڡ?ǥ�d4���w#�����y��1�q�ݲ�-�S����l����4����9�V�o���Ŗ�%�& 3��O�5��w�hIy3��3͌���4�6N��{q9�7��=�Ю��u��ޝؓX-�o��'�_��Ʃ�qZ��H?3���薝#����V�a<W~��_Q��(ܸ���N('�����t�N��b��"��a����{�8�{�S�F�KhA����I8��Ev��V��xÌ@�q̓��o�H�6o�R?���.K棝�Y�9���43�i&�3ݴ���~��ߠ{~C�	�G��#�,�0JS�+��EpM�����0-��s�Gj��3^�=N:�kAG;0�ā<Q6���3��;9=���w�}��S��|��V "�� �[3�!a��&������=��m�fƍ~2,M����_����c�A�_�0� �]����������In��v�{ �&IE�!ːiG���"�2��Rg���F?��=~�i�g�%^v�2�::�t�]��f�דw��ά7�d���~���+k������][�`�r�
��vc�o�9�D�sߢr-2��� �"���	��0 Lҽg�n�H�8��A^��@hKy�o�밙W��w������e����g1�F��i��|ҭ�3N��N7�x�D�˷<�O~����_���y>�������6M���m�>�hX�ͭe�/��R ���o��,��[5�繁��}"�!�a��S1�vff�7]*uq��*��V��d#sT�%bg�Q�ġ�Z�N�!,)H�|�6���'#µ�v���u��}��/�&�t��L3˞��u9�{�?��|�Idlᓰ�8i��.(oG��;M/�<ZO��oq����.���"��t=�L�!0�_|q�2j���p~��'NMNL�ܾ?;7�[�A����d��
���nT����:=8�6D��T'�O;����d����ie�f�t��A;��ݰƷ��������fx�A��6����f�,����a�.�;^��K'GH�5�uI��-¶R��iK�J��S�=˯�q4q��˗C�D7ÑO��g��g�ǀ96�^���8�iT��R�%��cۛ["����H�X�@��2�X�u�1#�f>R��v�eH�gڲZ�r7��mD�!?uX���7�,������6����t>P���ii�̇�9�\ƣ0QE��巔9��FTe5�4�OR{�VD��tK_Ǎ� :Ú�&Jӳ��#��Dt�9>~j����G"���Q�C~�d����P.U�����o�MLm�r��9o��P&�������J��#'�D�
�[ �0��[��_6����&��6�,�ț�~k���A�<ـ~��1}��|�]��X����I���OiSZ�h�?P$}Y͂x�oy2/�����y������]9|�P���e\M���<(��+�&��c�l��p�X.ӊ�X�./�5n��.��E�%�w���������햍����?Ǧ�Ԉ] D�u��!d���qoทh
P�<�(��T�TZ���U�����W��_do�p H��i�/.}�g�mxJ�Ko0��ʐ����D�U�ֽ ���".˘��K�gx�f�?ː߇��yfd;�>ᇝi�ݖU�����i�S8�c���e�8D��N۴ヷ�Ep��歟����2��>6r#��S���x;�<6��M]��Np^��)��)�`Q�f�WX����A���z���DP� ��� ��A�u<�3�t��=dh��8Y��/]�M��'h�$�@�#~]��;����01F
���t}w�2LFd�d��W��-S�7�M;�%d�]6_�S�H��x�W�Ɇ�ϥ������.:���C��3���].S,HvY��rF��P>"d�K�"J�SF��AjS*��u����T�4|䏏���`���2\�#�3d�V����2e���ƫ��ib�}|�?�@ϸ�^�#�z�F<M�1�D��3T?ƕM�چ�%��h�^
�-s8�g[��_��R�0?({>~˺��k��rmm�c�����t�9>rsF T�;�F<�w�߹z�����X������De������l�D^�&a�v�m���%l�Q�K�/K��6N	[�����)��?����K���o�W+�m�,g�d"^��6qL�������o�M�Y)��d*fݨQ
��&���@H���8-�5n�G;�Ԅ0�ގ<b]�׾ѐ��5�H���لrd�H�Ȟ,.������	q�%�I������C�IA2�k)�������ٵ����+U����0����zŲ�Q��!,�����u�`�H��P5������@���42�v�>��q3�ߙv�ND����&��IEu�"N�L�ș�l��_I��-�A֩��|hĤ��*D��vVM�e�O�b��}?Y�,?��I�L�T��J�,�0x�7�z;��u�v ��@s�֭��ӳ�o��Gzf�a6sHq3N��5�\��qj�\a�+�t3�Ҋ��T!:�3s+�4TVZ�6鮛<7�0ݾ����4�=����������l�3-��hg�}���M�s4����Y�^z�G
�C�*Z�!ad�|7X]'%#��w�*��k��r����\�(��3�n	�˗/�q��Ery�3g��fKN����Ǧ�c�{���b����o����Kw�./�z������fc��Ie���R�,�4� �Ү�{�~�[Z�}�L��f�A�H�u׿��<:�a4���s����w��-"��v���j��C�j:t\mөM~�~	K���#-`�H�q2������"��uGY?��-3�}v����g7ⷡ{~m���w��w)��0��p�a]�/��/4W��aܳi�VW���D��p���ͱ����nq�����?���~��G��_���%�,�xyǁ<����*^��a�he� &�cx�]_��%���W������ ��,Wc���P�D� : rn���I';D[ j\��Y3aB�,�s�D���R��f�.A��e4>�"D�eE��R,�\&��x��	�mo�f�dC�g���ˍg�����	�b*�
�4�4GX`��A �N<H������W�� ��n'�p>y����(�G^�W
#T"s�>�O�@h������RG�R7�i�4��~�R�4^|p�扽��щ���0u!�w��X����]5����޽{���8��}�'yD+���������;��O`�i�/`5�x+���H�:G�Ѱ�N��+�Ӯ��M�	�wʑ�Y�ϲi;�v�n��Y�}�ʶ�?G6�2\)���l��)<{�>4v�o<�a�?�,_�~�a���a����=3L�~�V�~���0�G�gx�&KKKA�� ۸�4���M����#��ʠ\���3���\������A�&Y�^��ʻ����~�f�0+0�,,�!X�`�
��bC
i� $�Z���/��Eb�3�XzLO�L���-�rz��ߩzo���� �}����y�ɓ'O��Pu34x �L"TXQk�߻���5͎���#��ߒwL�$H�`�.�x�E����o���ʉ_���`9vފ��۬�DL4��X\�]&j���D�d�>��s�%����v���
8i�#��6u�q�Ӽ��p���ģb��Nެs�_p������|l�;n�e	K����i:����+�m�󷣻0�	�፧�k������T�{��M�� aS��c���}C���m�[�me�9P ���ޫA�u(�� H�)��'Ț Ͱ̿�m��qC|�9�n������ST*� �'�:�yQC*W���{`���89	��	��!�\ۜeґĖ�Ɏ�&���AÅi:�$R���    IDATz2�vQ/kk�P�(~\:��߆��EF�"��n�7�#n�O�7<g��oې��?�1L=wҏ��<�Qka�ߦ���7q�l/��>�&7+��ܡ���S�o�C�
�>*t+p*�%\��@Pb�w��!��iZ 9@ƿW�Z����P���x	e{�Y_�,�'��[F3���~�%�Pm�{��y9W�v.9�:)p�D9U����(�6!l�Q9�Sۦ�G�-�Z�KyN���j�j�B$EK��N�����Z]�1�i `���m�E>�Ƚu�%Hb�q�V�k���i�!�5�_8�����e�[{��o���0�ۦ�U�
�3�7J�M��76̌:n�����FG�6�  �#�f���qr�'; ɢlP4>=x�˯?�͸��K?�I���f���2,�R�5�tƱlo+ST�N6k��v�q�[˴_W�hsnwNE6]�Q��Xyӄ�Q��<�P��5�Z.0�3.��SG�����00�I�n�lk�}/�j�*�eX3��2M�3N3�f�2���WK;Ju�R�m�E�����qk,�s[s��V;�~�(Cx����Jg#�a�9u�����lp��Ώ�>R������Ęqrk	�щ����!u<�y�1�O��wn��Pc*��w�+����Ǫ�@�Ͻ��e�Cekr@��`��D��Y���e�9�%��!acT&�d�z3g�trx5V��~�3^�H���g�n<ȸ|�T���n>�4�t�6�ȷ7FJ~���c��Lo�$l;�D�O�6���v�p�%w���/����n�_�At�K W�����M�I��?ٰ��6<1��4��;�3�j�(_��n��������-����׶3��29Zpb��1�5�#՟���N�=Y�?i1.��].G*+����!���O<W_E�����r�b-�J@I�v���8I�����('�ǯ����r��\l'��Єg���g�a�m��M8�d�(�8�.����~�4��Ҁ���靃({[�b�߈pX�m�o����Y�ܖ�����?�t�؉ٹ�Yv1T1E�XyS��_]V�J�x	�l�a�峍���3N�D�@�pަI@gj�!�s6��oE���t�k���b>!�P��E�qɸ�7*�������~���/y�;ʙS'�[�r��yzv�����Y��@T�O����g~�_��7��a���M�P�,��n�G���h��o��!���O��0�j��/jh�;@���y�j�5o��EZe)]ԧ��߰�'���y���QRF�O�L���V��h]��-#ܶ�0?yة��[��[F��z�_&Q�}hKX��s�f�gʥK��&g&O��j �ȡ1>: �uM��8�g<��7�n�����_$|!NB�� T�@�1qR�0��.D8p�]������#,�,/�I6ʻ�����|gy�����F�=���A\�f�7р�H���n��ɢ�n��Un����������/�ŏ��ÃC���7ʇ>h�)�W�];Kg����m��Ω(C쀭�&<~���o�����4��m�$Ќ��ɷ����;4�q�i-#�}�Kt��Uƈ��Y��ǟ}7[aڬRm-R� 㤳����O�M���È�@�{��g����������S�P�Վ!�3>P�a�	����9���4���c�@ME���㮬,w&4-n�],�������a�������3g�F��;������t���Ъ%AL�Z/�+Kс�ۨ�P��n�@�̗>U�㻾���o����� � ���#߸G�vKW����au��m!Ǉ�����f��ſ�ᨶ������e�q�m$����5��6]0�x�N\>F�L:��q�dX�M�d��D,A�F���x�@_�@{re�3�xß}7�!��t�{p�Ņ��Y�=������К�͜��I'	 l��?�N���̣Ǹ��N��n4�yBt0�^�hSG�8-v�&�,©����ʷ������?/���x��ܭr��edt���=�텐�Gǆ�2HPk�ۏN{��^��^,m�#��gv~�0�5������|�,΁L��H9�O�˶�	�KOo�t���:�Ǫq���F�He%����� ���[M�"�R�O��~�8M��	� P��6��f�13��X��ۺ��������3o�c>�x�˚Ag㼑`�웸U2o��ͱ����S���.]�|�����@T�Q����h�g:��8��ЩJ@����j琯�6���R.5L��w�ÕZ�u�G?2v�d�!qjz�<:V~�����)O<�tp��7����H�mM�P�����Kޜ���\j)�ss�29�k
��7�5���|��`5�P)s� X���A��o� � ެC���.�;�sQ�
\��=���6���X�
�J�D�m����a�*�/�z���:�6c���-F��9�tF^)R���0��d;���\Gn�D�ށ�m�d�Y��o�6'
��,�щ���-��s�6�����Z'^YjT������26"]�gC�?߻�6�3����8	@�ã#\?����g�BY�+r�U�?�ߖ�]�QN�8VZ�}{�vi��0�0�K�V�a�ٰ�_(�䱶��|�P������ksL {�3��.R��/����\Y�X(0� |����2�\F��n�3���G)s+(f�DR.�dm�KN�K��n£����L�y���4��n�_~�G>7t��诬��E�)�����D�:<dO�o�V�`�����'�li�966�+[V ��a$��?6��0g����{�7��"O=q�n~��Ov�9�=9�0����|��{��<������-�mO<^nܺNf=eim��,VʁC�M$ N�,K�a�Ņ��K�(tn�[Y[(K���Y����UeN:bIԍ��2�����C�-��(�T�C�O=���V,��j�=5����U�Xu�f�颭�X%��7�%����;Z������:���¹�o]���|�=�UV�6���89�J�T���F����W��{n~�d�}:�p�9�z��Iy��-f�}KK�C�����:�A�Z�d6���iX9�9��Xc�L�O���ٔ��{�,O��K��dp�<8Q��뾮��/�<��G���g�0�v��,hJL;=WO�w��6���ѰeĔ����؊&+�p}k�q�hKBd�x^ڵ��qtx�\�~���^,��?�n�zQA�]�ss�,a
{���r���N�=S�H�� "Oߌm�vO�)`[�.`%<������?k"$�vǈ|:�)v4�J�%��iį.�,�wı}�/�ŏ�0vt��2=3]&����9��훸�v���n�i��GZ;42�422�b���BD %"�UW�X��y�٨�/|�;�6y�="�'�bz�6��.��:9�����ȷ�3�;�-���o��������������-?�3��,b�8��X� ��eF��!؇ö�K�=�\�|�}�K+�c7������Pk�](]}��@��� K�uu��i�Q�G0{EDi�_�n[e�`wz��8p�<��g�����K��G?�2wg	9��ϔ2��0~`��۩6�Y��.m��+�.,Y�#����n��� M�&bL����o�ո��$�:�1L���HO��h|7�PW9���O�f4#��#A�L�[�-�����RYX\ w�V���ӲN.O���M����H�nB4��f�jn߹Ӻ35}�ƍ��rC+r/�� ���fx�U ��o��Wxm�������p�$�*/ S_*�O"�_���]�*_�~��'�SSwB[6�X�4 �A\���OȡoܜD.$��M:�~�et��������#�aq�E�ۓUMj��6S�5F��h��p9��q./��[�7^���O�x����R����-�{���0�.�=r��KmW���.᫖�F��$NF��2��h3����w�%<+�Ubn��;␮7sI��̞B��S|����5?q�S���1D�eĿ���-\e`��훸=f���2����JЃ�]#�肆�v��o�Gm�@�����{��ߘV����,�I�����|L��&��u��ˋ��������Q~���Us3�����7�!�jiK$r
��B�=��$���opS�2��YB�1��-#��b��Vy�«�7��[7��;�b�I����cTa�����9D�6��V1f�A�(;�F��0������ղ�:�:�U��-�*O<�X�uy�������k�X�Dg6V��c����d����
c���C��ֶ�D�7�Bh�1���vʻD�N���1$�T,��U;��Tg��ša�j673#�p\X�Z��T��"���M�� �1�a��X�`p�P>0q`��x"=�F�ƭ��׎s�`<�Kx�W6�����ɶl��^�t���2���P)���G�G�?�����_�;0Y�2�0
�WK����y�g��z�.�0s��M��S�����r����g�`���j��A�GN+g>����zp�"2�P\��*Q�W��[�f�p���z���/�wXb"�B]��Ï���vy�3/R�Fy�˞(�=|��?���eq���m�
m�� #��=ȩNb-��C��X!:쿙K���?q��t�߻�3V3O񞋌���nA�Ue�$甌Eݧ����R|:�;{߉�eD��ܛ�n�T��׹.Qi+nQ�S�d��eG��"�w�P�m`d��x�c��)�����5�~�cE�w/�2� �����d��gx������?�? f�@��Qg�͋9�u4#/��b9u��;dr�&����1uy�u�Y+g�?!v����˅K��(�O.�xf3Z��c�)�G�����2�`z��5��AȜ�;`��i'<|�H9x� ��iĊR.�|s�Vy���Pa.�˯�/�#c����������}���⫗�X�̈́a���KBU&L��qx�/ A�w=����t�:V#�s�?�m>Y�6����iS���$�N��By��-DV�;W������ު�웸X�:�����/�e����X�7�l�oh��B�S�t�5N ���ݶ�̼���G�SV�!�"�f��o��o.?�/�r���a]q������/?V�#O<B��GE�9oay5�mD��r�ܩ�>��Ǣ�}h�z��2<1T�f�ʵ;�����L�0�Va� ��"dx8uϘ�౔�v3�숽ě`Yd����-�
��a���4��b���+/����+o��'ʍk7�s/|�|�S_�X�E���/�Ͻ�j�7��
QJbvBg/'ﺀ+p��Y���[�k��F'yg~7��<��bĕF����S�ڕ�exd ����o�N��܍�����}7�ބ��J9�;̳S���.��u'��w���-� 8��O�]�3��qI.���څ�P*`�_#8�.�a��y��5�������-?�S�c9}�L�]���/UKw�߄p�˷~�{���$\e	�y�ܞ�Ew�����O
���W�^-c��T-��*C��f�E!���xU�ܕ	%�a��D�b�Z�Ů������ˍ��W4��3���s��XC�^@C32�.~1g�0��r������k����˷�?*���(]��_��/ï�p��MD�U�(�rw7��*�T;\Z�U"6<ݽ1��ɰL~d��M��ծ��l嶱
�@Z#�7��p^�=�&j����o���m�u�:+g,��ғ&�*ہD\i�
�X�%�jl���w�w Jw2i��8��W>�������1;����So��������Ν�ஊ+��.O��_+�,��6cf��<R�_z�|�._��_ZN�=�n�r��Zƒ����X?�ݴ`gҶ$:�256*m���+�s[S����W/�R�#b<x�zpN�A�d	�����X�^�a�}��Ce��hy��G��+����}ٺ]y������WED]߂q�F���>������X��I�:j�n9z^	cGфa��w �?�I|���m��;�o<�����̟��(�7�k��˪��ʚUP���/��6��Z��)�"	����l��y��WƬ�ĩX���� ��-�͆[�Z������[c^�E~��t�ޙ�]�?�H�ٟ�9v�� b`>	\e�ThZ��uџB�mT|�Ja�ň�z�tY�/>�e
N��?��+�g�8P��h([� �8�4;U�f�Y�\@��}>;��b�s۶�v4�:t�@���̡j��Q�Ⅸ3\����1�tN��[��}��K��.^//��jy��g�[������gXI=T>��O2�`'s{��y{��-����t�G�#�쌎����a�)q��I?���[���u�|�g���M�>DA��<MWEv+������������=�~��{A�p���k�*6+�j��k���+�	���֤k� ��d�K���۷��%L B_.g��aLy�o9��YA��s?����w��!m>�˹�t�o#W�e=�E.���_(G���G�-��w��/}�Xyۃ��o��8�(I�a���e}���$
6F�~�w�GЉ�$ƦD�nԌ�c�Ľg��5�Zc.��?:!b�,FC���e|x<��r���#��&-/~����|�|�}e9���2s{�P�o��o*�G���~��R���PAv��w��a]q �	7��O���N�8#��:�}$d]�[G����b�:0`+Yı�۷�o΀���.B��7D�KU��d	�sL����B^db��r/�  ��p3��s�L�| f.����I`{ԣ����1쒧r�:6���� �����/��������{�ɐ[����L;��=qd���xp���-�k�A�}��b5t����d�B��;��q#G�չ����$�z
���t��Q�z�\���jR�Ս���[pDH$d��6an_��m���i������c|��Վ,-!����Ĵuji�ej�/�_R.�r���G?X�|����S��O~�S�U��Uϔ?��?�6C-�փz�Is���Ĩ�p��ĭ_f�?Zx�G[�h2N�#�#.�Y@��������[�$۲�TN"�A�>6::�r�F��Hq�?�&n6�`������O�b����L(?��c�r�>I�����!>�����@�u���L�o�3�^���Պ���0;�����?F�mv{��L,���E�$�~G��ߚ���x觗]���?�ɏ K��'Y49|�@�'��׮�ZΣ��B����h:�Zȥ=|G⎉2V���D�	�
��Tn�Q�:���T�F�t�W�C3`۴� �5��W!�j\�8x�H�9}��_%���G�'���v�|�g��o�j��+���[~�W~����kl��d`n��U�J�6��u�Z�^��vV����7���o��_~'�7��;�x��0�W�b��b�żzt��	�n��=҉�S[ �" +�۳�aL�P=���q	 �l���#˩u�'����_�k~�|���N����k�c�OS���,����Q����I�\�}��[AE�_dw���#e�=SfYJ�ӟ.g:G--f��3�0�2�tKM��0�V�vG�L�Xu�@�j�f�PB���E�=t2H��U]7D��5aD�m;�E]{����z���՛�ባ�ߔu}��By�'�j��+�˥[��S_�ty��"�L�Ǟz�L�b|����u]�đP�x:�Z�V���Q>J���:F<�4q�'d�w5N�%��ȗ��v$�q���/��'9�D���k�9������[\��o�^n�7U�"�޺y+��yn/^���>1b�3r�g������o��t���w'��oôs���lC��
_pRc���7?���=��&v�L`x�b������7��FO3+!_�6#����it���aӱ�A�,�}s�:K����Ct$�g�<
D�K���d$aS��"R�7ce>�!\�Y���4��h��1;��h�cP�ҋ͈�wX=�0���{ј�o���g�8Sg��	?�Fe�<�����#�ș���W^/��,�=��5�[�X�D���?��r��l��	�čL��u�W	N&�V\    IDAT�5�6�Q�.��m�fX����;eV%@�;g���˗#^�/ 3Eq��p�pwS�w������\�p��%+t�����/z{칷�I�6R���x�w?�0�����_~����0���-@��D��?�c��qrj2��89GP�V�я�fQ�E!h���?�C�Ҟr��1�Z(w�$��r��A�#,��D|9x�P醐{GF�h^*�;FG&�ɓg!^�*�:#�;���\�[�a�{��G/�^������},"m"֬l����$WRG �^��[,r��&Y�Y�.e��>��'��s.�u��W_cԂ����uy拟.GQ}R�O�Px�q�.��q�c�B?���;:�,��W��N���V9z�(�EN^��/qc�?�C'�7����7F���g?�kiq4ڞN���\���#nd��A�lN�+�;���4i�|"��������-Ӹ+��~��2t���V`q��I���Q��}��˷Xf�x����g�!��X��d�\�q�̈�bM���G@\l&�hx)�S���hvy�6jŀ���E	C��K�۶�"$�.Dq��X�uH�� ��01�\ԛ$��!������X�y�v�ڭ�V�5aPn1�@?~��!�$��#���Yn_��_U._�T.�!���&���o��7�g<ã=��t�#]�J|�<	%NƋ| F���T�:E�d����B,��ٴ��+3��YT���g����Z�*���u�!�Ǭv����r��;7[�[	eE	@B�Qx���r����$�rFc����� �+������ �mZj:�?��B��;W�����2���Y��W�m�%�vn"�ݙ�]&O`�U�7��?W��6�c_�X��Q���e��]6lI�c�^�w!E�E?n�\i��6:f�����Uİ�C�?N�<"^L")�{�:��l���8�~���:�?�mN��S���#�SNkh�^���EwD��0�]���<�m����O�-�?�jy��Ǣ/������>\.��>�N���d5���p�zhgM1�&����#���c�S�m��4pD���G�w>�|�I��㝂6�p�g�OcW�[}23���c/��!n�cо��/qo��3����N�!P*��v�>���h����x=4��S��߫nٻk�#�W��۞/ �ܷ��&�9����uo�6պ�)�����(7��pX΍����h�����by��M6,�DgfC��u�x8)5�6D�2�\f�c/m�u�����R��3�l	T� �b�Z�,��a�����26Z;>\
z��ʜ���H�7�!g֕M:���vC5g�l��WY���|ײ�0���s�4���S�~�Xz��'Y�����0;�PR��a4H�1� (���	{�xI�gr^�����q���㛯����3/�\��"©�y���,���X�][�A)jX�#G��[�o�k �����t���[�l��l`>��o�R���@nz����\y��u:���'d}��锹gf���6�Ͻ�\y�[L�yЉO�Yw�?y�:z�u����6�]H!Zx���7���Sw�%�E�ι<h%P�u#���mq��ۦ�׽�N�5�b�[[�艇, S��c)XB���g�0sa�sw���*���F���~�3&���7nÙQM>����/>W�����(���-o������ ���%�L���n�$>�đ��N���t7��wtWI��Y��������%p�7��f���/���]0D�n !8e!r\��>�����Y���A��葮H���a>�݁c��{w���4WN$�y��?��1�΂��� �E������ٍ��r��q|�\�v�vk5�-ƙΔnV��[;<kw-׆W��axU�F$�Sk�d��VUY��w��]C�-��~�#~��
c�oa3�}�ڑW�A�����!Z�9^ �l���̅!��FY]� 
},���"������?t��ȞNl�~�����ʱ#tX����a�_x�,#�n9v��:7J�'��x��,wkP2�n<ݝί꤁��q;]0�z3�LI7�0��`�V3i5�[r�}7̢zƞeo��67��>����Y�$���H��Vmf%���[@e�0��7"��c�ݡ��}�� l{���c�c�6G�D�Z�M�sp����E������W��Ȳ9m���n�m�8�V����О���
OèM�z�,t��J����Cs��݇ȱj$MV��w�j�$�i<�P�B;W���.�ۑ���@n���!p�U/��]QN��v!�r|c��W;����=p���U^�z�<p�2�>�.gΝ)/>�
p���.q�L�^��w��q�2xԏt�eG�%n�u(P��x��X
�v�&̛���8��� ��V����`�CSiD�&r��lx����-�i�f�ɰ�6���ÕFw��)�W�D]l����! 츽K��6.��v'�g�2l_G�
\}���D�]I7�,�s!(6 �Hp����.Z}��Y^nn�`�ǈ�[M���S��'�Jؚ�
�8�U��Yͅ�d��=�
�|�����ܱ1��~h;89�Ot���тY!*�W(YWG�뷯���0�������?�YT�'����?�hy���uz�2���`OHGb�9;p��(D�S���H�������0]�c�3m��N<��ϑ݉��u�rY|ۦ�f�o�:`x�Xo��"�8�G.)wH�0�h��٘l���>�	Wߦ_5ߑJ�G��f_���|��} T 	�:�\Ἶe8�;cf�/_�T>�z=��<�!��!��%���&���e&|څT��#R�c0"'��p�t�y�ܶ�Q��<�xp�?^F��YJg`�G�uT��>�B�tT5-��:�|�!��i�o~#�@ �w�ࢢ��v\.��C���6w��E�+}���qt����:o�j�l�]��h{��� #�b�6d&��th�r��"d��|�&���?���0��3�;o�+�G:��,l�.�<�;a�{�Ľ5>�օ9�G�HU�>{�lp	�J�VT��I���ݰ�w�4��yd���%}�;�*N\u3�gjP�����nZ�V7%�m��+7/ý��Q-(�o1�rgMplf��A���JH���q�25�A�ѷ�q^q!�4���=,ǐy��4��6Z�iF�ؒ_���"C��^B4�*�ؽ�́?����+������?�8���7&�pl��HΈC��I�ѻ1�y�P/։�L��f&cdz�	�G­xPmWc����8�@Bd
w;�m��4�M�\G��1މ?�~���<���w�'��`N7n�(ׯ_�<�0m����֤M�Nw3��~��Ĳ�:���6�G��_�5_"����a�����l@�ec}g\�(��g޾M�oӛ��l�yNc�t�/���"�+;4�EC��>ȉ��h\	�=ѻ"�%�"�ݦ��/bҪ�����D
�3�4xB}�\m27:R���A�X>zQ�ͳ���(ps�N������,�ϗe&zn4�]��7�Nx�\���\#��ɽa�n�v��x��v�∓N���qք+pp��8�l(�n��,@qM�.'��{��r,�,���@9�~MՈ�OpjzM2(�(�+L+!JĆ��čp3N�ķaMB׿�.���r|�0+N�\��o�kq�'��Mܾ�{dd����JX�C� pO���$D`���� �1�$N���o�y���Y9L�f�D�q�?:ĮA�'E�(nܐ���{Y�^�xV�!�qs�c)g�CE�ї�3�`O����zƙ��c��Ǆ2���ȔWm���pkb|{k�D��Ԋ�n\��o�;�e���[lfq�>��V*>m�
���/W��W���s�F���U���n�	�~��aeՑ�c.^�j?��N�+����g���2�<�����A
�g�w�@q3�/����@ša�G��4]������m{9q,�:u�T���{i�c��j���9����z�������+fu�*���0%��}��Qy�6�FAST�Y}�f+�8�q�O��?�w �]�r�U4��4��TF�)�&�r� L�9�A���������tp��FP+�R���P��^ۼ�������7V�'����y��B�j)���W��[#�qW���.a�@Ⱥn��J����AڸH��Ȋ�ת0t��o'���K��l��r/b�O����w�	��)�8���q���\�!�	&�m���<&�k�Kݿ#��*�����r��U��N<�����������y�o'�jJ\\�a�8����\�|o��K��?��	A���}c}��	E�V\�'����9[Q������&�鯘��cK����	�R���y��7~�7F\'fZ�b[��Y74x����Јx �;h���%u-����ۊ�W�U���2��gr�(rl�x |yq�+hK}�n���y�bF���ys.�*"��q���M�Uֹ;`$����?�g�8uJ�S�{#sR^���4|��4u�j�7��G���+�ۮ��Ƹ��fp�I��y�|���娊���8��5 a�?2���1G��y���y+׌�� P[���3N�Ź����:�S:��p6:�/��s{�#��A[��pP�w�F�ج�o��ț=׼m���trg��v��3�~�y�~?��?�&�r��T��c\ۆ�8D��]PT�c%���fPNh'��Ғ�1�+Vݳ8��"����������*>*�ɟ�I$P�Ze"��i�'��lr�D�N�ـ�	)k=�YU�M�u��Q�l�v�Q��<�r����HG�u���$J�u܍�h��q�͵'Y��V�v�q�Ѓln���	�g��=|XUj�E�N�n0��¾�$��'��ﬣ�L��淿���xQ�I��n��s���n��#�� en�ەH� �;w.& %V(�+���ƷWJ|>��Cg��w>~擝i����8Z�2�zw�(Y��Z�T�\5'KL��#�0��H�dzp��,�q&6��P!����I�N��&MZ���Z�8�n�Jc����R��M�/v��:r�\���p^�#��i��m_�Q�\]QMXȤ�A�U|����Ś��C9w2ML7�f�G�!����q��.�{�n�x����ʴ�ru�M\�N(�����,]�:����?��<�-�ģ8�F�W'N�W�YY9�'q�W,	��{�u~�=NK��iNG:�p��Hl���P��F�[i+o>w�7��Q:�����mfNN�F�4z�ɤN@̡�0m�Jױـ�(�NH�[���RX�!bH\N���ejy�^L���L�B�*���N��@�=e!;�!K����|X���à�3��Lԝ3�T����-�I$�@��� `^�e������ꤒX�W��"�"�(/�����­w���z����3�Y)�=[����Z7�x�z�>|s�Q�Y��Gv�0��xO:˭e���������^��ү���_����_|8��c�$Y������so(s�����X	���y��`1�&qZ)�~f�[ �[?�C��o��(��<-[?˲�ۡ���1���l�8"ӎb����V.7�"�i�N�\Sa�d��O�S�b���y�rtȝrn�M��z�5S���ud@�ww�
O�S����@�:����/��w����\����E����aX�9��QW���>N��n�]�2X�{�$H�`'1^��cY�7n�e=�m]~�n�l��q�[�ąODʼ���z��g+�k&n��/qCT��=��+ �E58�N-q���:Z��z��)4�I�@[a'8"N�	|+l��=T=��~"���G�F�-|���f��,�Y���*�}7Co7'��[f�N�����nsvv�{�	ey�O�b	_]�`����u����6���#����G�*��?Z�Cp4�L�>��P[ro��͞�����"g�wqb�&�1�g�B���M����e�	���o%2`����A�5���vb�(&���ݎ*t:�2���ު��B�k'S����g�b s���w�GM�@}5,S���/�c�+�k�aֺ*G�]�`�1�-�"N`!>��Aa�u���l�����8�m<�|�ʫy��+3�m1��p7Y�P��5_�n�a����;	�k�8o��K�QqKN�!�H �>}:z��)FH���f/mt�SbO��~�%�$~�q��ϕ�U�\�>`y�V��.����\N�,�R+����'��7���se�x./ /[?�thR�Gʦ�%�;_�v�{�E�И�?���x�?]��A��뗣���Qb�D��f��z�͵�Ç9��)R�i<�1��-WƔ��e�����eX�ɷaͧɸ�o�.���ā�^���辐KV�K�Q�GU]�d=��H@Y�l�a�����<����	��ph���&׶�Vݰ�D��䁚�# D���3��.o+�:s21g8^�Su�+��������G_<ZEқ�h�y��n��.��Ṳk�!` 'KgX����3~�;��rP&��(y���]�(�y��+�^deG��N_�92���d��K<>�ϝO�~xêz����m&m�E�p~q-���0d����y+������}���E&�[]�2�D�+��R�\����S.gX:�� ʷ��	x�D�.���;���VW��"�H�ޭ~���,u�M����g9n8Xw�(a�Ѣ� @��{<�b�5��b�&�t�\�6L"�5�zA�Q�=�ؖlF?>���m+~A�ؙ&�u��l~7��mÞ�	3��y��n�D�@hgU1��&�Z��<��O�۰��o��x��w��v�^g�O�Ȉ�J��7o��u�4����CA�
��occ�k����܃�m�Z�X"a:���V<���o�.�ˆF��aX	T�'�;[WÀ��f��#�s�w/gs��42G5$�&r3`�p�|2�A�ڊ���"W,��rc�F�v�R���S����R� 	�oN;.�HL�сb'�F������>FM�*ڪ8$��D�-;Dc�S�c����D�;��>�%l�.�!vۤ��Q,�yZT��L���8��w*,�m?�Lox���������E5�?�$�[gq���S����^�
�{�|~X��KX)�Z�"B6��It6�	lM���8	�f��'�1<�c:;�gS�>�9�:�f��$�-��b7��� nI���)��H#�-�eN�0$A�Fs�N�S�\��9�\�O⋣�E '���{o�[�!Ĝ�R�����v]��w�0k��l�)���W���D��^�M���Y�FW	��2�ϲ�S��Y�5�߸鯟�ű�r�����/�\��IA����&xwo(�I�wP����o�c���D�E+?�L];�l��|��~� ��H��wܐE<�~�o��GU|:;�y&p��m�vܞ]�VŹ�����B�ƸA���w��B�#�ߛgٚ3˥+���{vӭ��h趰�Hul�u�o�=���(�<L�B����M'R�o2śq�pk���ٮ�.��M�c Nʹ�U�~w)����M��w:��N���?��۸Q�J�y��0���6���#������K��~K�)��s)\��^Ugeu�;��^����|���  �K`�n"�o��!V��5���tTB���f�26;;���7�-��$j��˵���Ԍ���._|���q+Xj_�6����кHt��؎h/�t�M ���	kM��#��6]�G���t�j&.5ϝ��"y).9Q�d+��S2��Q&d�M|BcB�_�3jM�IPg�a}��䍸Q�[�i���v` ��;
�ߑy*UF�u#ORo�Zܥ�W�>v��'Y1��yf4s��������/�8޹�H}�9��<�z��>����:�[��I����� ������Z1���ɫe��+�`♧H�\ì������[�٥�ȗ�9ْ�E���V]=��fh`\���V��i�>Q9�@��m���T���$���    IDAT�"����ݕ/�ԲjyvFj�����3�n���t�[�D����%6?ce��Cq��*A�&βl�0�O�ee}2ܸ:�3ν�#R��L�x:w�\�H[�np�ihMjo�{��7q�����0�b���$UoVІ����a�K�>��۴�o����P߆�N�o��S� B@��<{��=��{��oZ{���q%�2�r��3�l'����u�'W��X'�Y7�u��t��p�-�'��L�w��v�$�����2?���B�pÎ�p�5	.�aF�2��pgQG1��^�|�/�U�f�(3PP��QF�%�������W�%2�2'���O��������7q�8�ծUO"M�{��)sأG��s[)+�pW�[D�X	�C �gw��&Adߵ�TM�6-ADi��v/�-�܍���v��S��)$��DU�79��H�WC��Nc�j�U$��q�G���(/�MK��H�[��55���!
UTO�Dr���h��1�w��ζC�~7;����8v{r�ۣ�U� �э���1ɚQ�_�"t�*a6�%Y�,�r����V}��$ئ_��|�Gɜ��ܪ��ѷ�M�u4���o�^\��(�C�	���/�D-a+s'w � �o�M��?	�8����Ir����␳j��n�r��+���k�D�ܵ���G��C:9v��1ALJ�Sw���QY�C����ݠ��YO�p0~�)��=�&�7;�u�~�����L+����s3�� ��vb�D��&N;��\��E4���
�if�Ik���wʾ�\kgX�1��w>����mJ����V�Z�Y)v:*G~&?��{��ƀ�~������_�P�������d�<��y��	�b�E�Kb�m�D��x��ƿ���U>�W��p��� !"_���6/Ü���e�,W���Q}�#�>��f��s���zsø��DE���E)�H���@fT����xUd�|L˓�Z��W-G¢^�����|��+ض�d|�ʡ�ġs��\���� A{є����p���&%�!�#����E�Ο,7:����i���1�D�w:q��̷�X��K'M�kGcӰf�>�~��C6���kH�v�H`��ʲw9|˥tV2��W����4�_��6,���@棿�+7��~����y���>=����U�7/���?��D�dS���qm��[��p	X�K:��+�'�y8��m��g;��v���!�ng;v��1���,+�Q�R�ɽ%p�77�E���r��Wr��?���f����[<6?tڴ��Y^�C������u��~7��ͷ\[KԊ��,�!��h%�f���=���S��(�W�M��%2�<��F�Vfˊ4ߙ�~"/��_��~"!�d�v���Mf�٣}�]5�ҙ^"�N$��[���o��+�FԈ�h��m�ۘp�屢���+��}&�RUM�,����������`h�rl-?�_������s�K��~��X/��-A�]�-�[��ϕW���Nr���Op ��\[!W7�OmCe���#-��?�����j���n�f���uζK�rleo��S�sc�Z5{�]�Y���*��j�d�Y��w�V8e��n�nW1��(���)����Ĭ��-W��4^e�#�V�{�ز�鎥�NW�u�[�,����=q6�)zYO�ȩ^	pv�3OãL���.�f�Y��w�hr�L��������,/�3o9��6���ܹs���[1J-1�t2��1^���M���N�e5����n�5ͽ�-O�[)�]m>�0�Z�Ú���;T���g7�b���.���_*/��*�a�,CC�/w4^;\�T��𽡂�6$A[7+-&�"�2�� �����K����v���3n�nۃg>��gم�7�8����K��#`Clkh����.�Or��&�؟�;�!$8��;�1����r~��s�l�8u9������K88��
�-�ԌE$�F���s�\<`��U\,aBL�`My���E���b8�\��hÃF�7u��c���\�D'N��� �}�U��]�p�a�v�-���(ko9F�=��R9�om����x�!���X�c�1x6v�{r����N{7)o 3��^�������1�|�g�~�ֺ��{	�I�,'�^s;g�p�U�7׻p�}[	Z&�5О��T���r��8x�����aE�N��X�r�2�k������I����	�㷆:�����L˰<{�K/��<1�ɵU	Z4�����M����	RYo��\[�S��H��>�qƣܻ\v�fź�f�ߺ���ٮm����B��m]2��|"���6��e[|r4���G�˷��0�-G����ə։�pS���6��䕗^�ޗaL�N�~ۮp��|u��0}�c[��ߝ��_�8z淿~���Xݶ���r�6�=�3ܓ~����B���D���_��awۼS�(&d'�2�B��ߍh�m\�v��#�Ry�2_����/��/���8	`��=�Wm��3��2p{;�� �E��;ʈ땜��z��w
�a�躇�X���?7{�k�	gi=K}lK����lN��u֥�}g�JX�q���|��R��[<���N$,�>5�e:1t/h=�MR���Q�y[⒬��/E��<�����N�td�"�c�C�GM��v�K��߸�O2ڍk������%n�P��`*�-�{O훸ٟ�α
}K�vEP��u�vk6Ԋ&��2�͸�N.p�F'�/�Ti��s�e���O~�\�u3��L<�X�������d�"����I�|:!���p�SRo,�t���{���#�7=j���){Kt�:�V��N���#��X��K�Pm�Y�z���]�6��0|n��_Hnz��x5����M=����]:�_l��N�W^y�56>#��+w�"��;eG��~3��t@�eܨC4h'e3<}Mo3,���0m�Th�=����2��.8�n�Ľ���Ĩ}59�e8t�w�}q��L���������x	�Ls�w�y�9��〕C̡��|����=� [�Z�fc������AҰ�`�T�D���x+'ֻ3Q/����0��T���\#�?�+���X4o �>����|���}���5�a�>�\�ݖ�a�����������h��Mp�J���q<���B>|�6�w��8�[�<C��#��y��� G��Wn�Gy�|���C*�@���H�ȗ.��B��'YՇ�&������%!�q�/��;��R�b�����A�*-EوB4���7q�goO���S9۞%�;	���o%0 Aq�)����Fuz��q�&���;�gy�^�I˕s��O�4G���H���V�>��߁����|Cq�R"ϕ� (&O��}{z��E08b�]�)�.��o�^�8*�KW���[ԩH��8	�k�$s��^,$�����x98t�Ӟ����f�� �ND��#��ƅ$T�mgKD7q�p�~ �+�߆!��;�+^�Eы%8��3Uf9�����}��0�]�c�7�R;�"���F#����������C�Y7�w�=������f;$b���y�����g���O�	T���n��7O�Y!�}�.C��+	׳��������9i>V>VOi���l`�8���z����v?�@X�Vgի삯r.܊�u�
��96ػK[�8e���&ǌ�,�jb��K�%4��j�Zը��B�X��ߘ���dM��o<S�s�u!8*�-�?	���QB���7\��	d�M�!(�@I�5pD`!l��`v��-�A�V��?d����/`�_F��h�J�:�=��o��Y[\/�7�b��ǅT�}�����O�K��+Ƞ�Ipz��Й�E�#��7�	{��k��u�����;��|d���z�37pB̂a�۶�J��-�l!w�W4�$w�}s��ծNq�V���F9��7��YBO.�\�4�o��N�V��is��pe�D��/��b������K�CTpqb�[\��� �fń�yVV9�b��� ;��zk�y�X����ҍ^����ٓ���4����y��1.gT1�~�J��
qu(̥�g=Ļ��1[\�4ȁ<r���4�^��1���G��V :�suןmx@d�Yj�7��
d0���u�������E�?^�\�È�*���[��[pm�	8x,���dN'�Vyx��}��i�8�#L�����u�����8Qu�v�����豣�(�A�m��Ia������}�t�ݾ���oqu�pͳ���ie������r�Z� ��~l`r��Z�m:�H��F��.{Ɖ:p]"�k:��P>��R�[�C���<������G9t��pc� FVc!����c�M{�@*��w����pu��Ŏu&��!������S�����8|�KNQ_��1D�@$Y�Q.`�Qmp��P�H�p��IJ��-MP٪C���$x�Nݳ��+��|�vh8��ryul�`�(�$pU���)��`�(&���F������ܩs��+��3��5�U�V,�a�67�
��.I��{��r�?�q�E҄aI�$��s���o��߰��Ω6h*��Fw��������7q�'mJ����o%PN7H�Н�ԙn%��K?�t'��o��rM'���=���|��s9~}�Vs��y�h
N=�PRx6�"|b�@��$$w�C�� ��,�I�A����9�n�v"9�?Z�:Z;�Xy����^�#e���>�l,�l.s���?y�s^���yp��yʀ�b���)[{�|v��M�Y�mN
1:�)�r$�ivr..~z���с���۸�ҝ��2���+�g��d9It���,;��Y�ߖ���+�v��y��v8wG�P��B����;�!;6S���q��[rY+i�V�ڻ|Rl�W���@ɸ��f��%P׹UL �2,>��������������rszZL�Tz��\�̑����d�u�n�lCn%����X�Ȓ�VBi2R�\1@d���uTpX�.�CAf������_�=��n"�om�Cd9��8-�1�ж�f�j�!tdQ��8w���!�)u.�O�+��[Q�.
9��Ӳj9L�7�ަ]T~�Un^�,�w�}�ϕ?���X8h�1(87�pw�\�C1�_�[*gV�Z�	�23q'>$8�������ɟ&������x�]��x^o�SIa���p�.����#]P����b����������nŒ�p�����mY��w0�;��Wy��M��D���I����?��?-W�ވM�n��PH�=��3��1���9�D�]����zH�I}Sh����!�3�X$��g���nq��틤�k�q��� �S�l˙�C7�I���ř�Y43�(���V���P'Q�N}ýu��rzURS�P]�b�"2U�F�7�ˑѣ��k����2�/��"`�+����S	�I���I'��H�h7>��W��t��o]�g����߻�(j���$��
b�����/qGk۫�ݷ�Fzjr*��@>� ���D�rm�����٨�w���Ȧ_��0ߙ^��2�� n�x��������@���Ա3�[�0�����ʑ!�jXG�B��d��|j�*�;&���!W������L'��]�нn��v���9Y>��w��xf�8�gl6F{�˹s��x�<~��r��s�����^��W�"WDQ$��A�l]��
��PE!�ho��{���w��a��q���`�~���p����;��eu� ��=�\��~4I�����WGa����
|*�Hx�7\�껉�꒸}gx�i���3�j^W����}sK��)�엸i���.��Oy��ڳ0֪ܔ��lP �C��N�M�/6Қ���
$���i�y�	J���~������D��W�T�a7��=r����Ѳ:��{���P�ü�~��&�P"d$�W�"�z�I���-c�����9��'k��f	i�z".p���>B~�r��q�Q�NZ:��J�y3gyj~BI� � �W�j_��W�Ӈ�:���w�O��x�|��ϕ+���:��n� ���ݶ*;��Kg��m���5B�8�$\�.��۰ģ�����X'��L�f���X�ż�������{��f����nz$�P�S	��m�#A�!�ފ��C\6��8�Hn��q����U�19�,�i�,D��j�1�?��?���W~�����XH���c9�ti�vq��w%wX{�Z7GE��-OA�Ր��B���å'XY��q^��o$�z-7�|���r���rmu����2���7f�x��N	��8¿r�%T���@��;vŬ�Sm[��E�bI&�Z�Q%D*Vc�l=���_�T^���+�����?U>���R�c���f�GV��Q�����m�"���$��$�H��G���o�mx:����.rɠ����t��:�2w?��J����1�{�=�HA���D�C�×C��3���6"9\x��?�������f�~�q�݌�yq�x˵>�|�	��~����o�	s+�y��������s�|(�^���в'�c�d���	�3�4�Ԡ����v���u��%u��u.�����/��bl
�K���433W�0����r�0��%A�z]rdvv���	U���������gQ��L͔���'������5�E�Cr�3j@ےb��ّ "�hu����K���e<���W�/�x��t�Z��X�	�7�
06;�g�7��͹�scas +CW�)�ݙ����p��;�n�Ww@�p��
_�/�t�A����G7�Э��2�ωc/�xx�z5چ1�3��9��|џ��(q����k�ч���6K����(�����G9�Z�D�6�[foqn���4� ���Q�@u������6�*���B�J����䊇�7��� ��u�2���MN+%����rm�R�m�pV�+P=�+ޑ݈p�h����Ux�����ӣ�f�,3�`1�=�^�/�˭����semv�����~M!��N@�4B'׆���*p��l�)�C3�RȰ|�E�l�SP!R�%�@"����Ы�6�@(�Ǡm&��������{�?��EW'�:;�� n��D���M�ׯ�o�>ӷl/?~�DؖhPW&Y���I�:��]	�^L�q�.�Ѵh�qu�O~�g�@�_��B���rQ��
�����8�����`�:9�8�e�9{r�v�u�v�89���v,�$�5�5;�.���)3��<!�Ц0�BcA��m1-HOi���s���@{�� R������-N�rG�m�^(���*t�k�9���enj��$��K]��n�W_<_Μ8[�������/B����֨1�C2�傰Hx�{w\�?>��ѷ⸎>�>���7Y�����9V��.(�����k1�t��a:[�;����{{�_��F�� ���'��1>�qژ���I���.@��~r[�ɩt�W�~W�.���\�NXݩbz�:1ar�U������+��e�~�B�<�2�|��������=�=�`�eD`�l�GG<{л/����M�£���`Yx��V_�N�k���Ӻr9��tX�EMm�Ё1bূ]�T���U\R��!'/�.����L�Go�o�������3�q�do������<#&���C��,�;i�~�t��&a'1f��~g���δ�[:G�A{lR�Q��3������G��8z1�o���M���#l���Tv�+*�99���M��`)k��h�qXAiu%ʬ�iz;��@|K$	 ��[�t	��9|Y?;�������{��ʅ�O��O��|�|����Ӈ���p��5�U�O_A-ȁ�twޯ��vږX>���[�R�S"���P��z�0����j����xD��Z	Z�n!���'�[�c��hUa�dvy$1slX��D�_�*7�~���w��$6�k}hHʟ���J����[�>f�fѐ�}��}��L+>�	�8�Ig���^�y�����/=v�"�i3ú�    IDAT �U���k�sit�f��E�Nό�7��7q��9*����=0\Ua�"�z�⎎5&[]E 8�����8�k�$��0�m�,���@�5� �@����ջȗ|�5�C ����st8��|=n-'�����_�u������ϣ޷f1�Ef?:v���2�Z�
X�� ��H�؞�N2��٭���v�7��[R����TL��G�:���/Y��%�A!h��c#�GG2k��1�1	��1��0s��ђP�k��8�Z)�_�\�����l�{�'s
:ê�C�[$��wϰ��	�k�a�'�2M����,�g���t��;:*E)�_��,�tҀ�]�5��v�|L�eV�C�l�ݛ��Mܫ�g�8�v@��ɕ�]��z�Jf�k��oSQ7�J�:+nc��6'�9�����o�3�N�z��(2�#��۫���3�~�)綎��^W��k���I�W��g�?Pƹ~�{$��<�h�=�-����5B�\*�=�,�l`qG=)|{�o F$E�Q�_�.T�Zo��h�f�����ǎP�4v�vR��͌-\}��E��l�;m�V���k�[,V=W���s��P��_��r����Ԃ8֗8��z/�]K탸rgRQK�0�w�~�~	_q�8���7��UmȎ�p��0���*T?���e;�vtpqI�J��[{�}���rWo��qnr��~�#)=�Py�W������:�买U q*j�A�' û6V���1,Uߵ��jK�=q�����{*��u�1q]���8�)�1�Xj\^^�ʼ�Q&�p�|�/��q������Q�X
*��'~ۏ��ZъL��dG:mV�RdmU@�#�ڛ��8w�BB��(���3�5*�o%^\[�5�י@�[t�5881bċ���h�	��j�*�`X6�z���Wb���ѳ�y�>���,M"�@��u��4� �0b4���)�#,�Pߞ�&��*��T�Է�ť��N�藿kN���9_�<2���Li���\���ҁ
	����#��#�8���o��M�1���B�@T�B匮 ~�ӟ�=�w���!����R��p��r�^䅿=4�@��	8�@'����N'��|�r��(��	�ᳳ��� �����G~�Gʷ|�{��M�e?ʦ�1�D���̵�r�vc��$�z�v k���F�h�	@]#��#�m5Xyny\�g[i�Wީ��@�|��Z;�Ҙa"�06>`����ȝ�˗����Z�.���W���>,7�7��>^ڳca��.x�Ս�a�a�2B�p�_x��~r�7L���~���S�y&���8�R[��<E��l�oEH�9��]��1�ƚާ��ea�t�o�~��?]}��^����'!}�W| 	��9����V�r �z�(�Z���I�� �hq�S�J��-_������S�
�r�� �E��c�t���Yn��I}������s�S�Ї>T���/��� r�Tg�f��'Cf_Z熭��r��58�������!�@X�ǗW�P�y��u�Um]�(KH+hX�]���u 'J=�x��υ#���jL�jh#��ln�D�k����Y)���	X����K��Ƶ����kat�˽�aC�]�ZtU�:G�g�8z.#r)
�b�ήq"QJx�'����6f�ڜD�针�	�����myvj;^&碘�^�vS����I�,G}w:ӢAi�1�60v��M���n���Y����3����~�޳O�ɾM !"�"���<ATP?}�y~�� *���""��""jD6�����ٓٷ������NuM&<qC|/3V�s��[�N�:u�)�*��@�f̘a x;�Gf^�L1���p��0��*S�*�@)Bj�_=��}2��5�� �@�>��x��pd�����m�s?��O݃�/߇��aG�V[�S�ftӛ�E����d���0٭k{�mm�*ca�����Z-����ڱ]�M�1��W�`[حl�c��k�������]���Q�&!���m�ZI8P��.ߪur_��yb������I�_Ӈ�;�l�k�`m�?IFB�$��aX��i lh�/B\�g��B�p�>}�b����p/��<Nm�lH��Ƞf�H�c�h�g\c�$#��1�X,H}��g����&�S���(ekY*	�aS =F�o���"�}(�^)Z�8�j5r w��ÿ/ @Q�O�eQBCC-�5��&�A��YS'��l����>[�{�J�|��h_w�.v�fN1�f��i���]�ZvS�dqS;�����۰Z���F2'Ys���%�B��T��nR� "�A��t��#:�X�qc�\^����lB�����w˖��e���n�ZQ/fb$x_��̞�p&��$|2�30�g�&ZA}����
ভi��j�жCi���C��7���jy��,^��V`��<`]q3�3c�,# �i8��H�1�Y����Vk���/ܬ��(�SӵЊ�}�Ī�@E���V*��b@ݹVi��7(iQd��M�J�l�J_����>6���K�c0�9
�����>>qƌ�V._��~��t�[Np?�lft2q}�6�DeЏ��aNGsÎlھQ����."�W���+���=����y\)�s?�q��b�䎢��ӭ\�B&`/��L�F���g�*Q�35՘hOL��q{9)~����� SE�o3G��N��6��B;���#<��q^��C<��e�%~צjM
Ħ޲O�n��p�W��
�	�ia�=�Jz"��WHH���H����:/_��-~�b�: 1���P�,篋�s�#����c�$]�Oh0�6��
fqD�U
?��Nު4�5.Ƹb;�N�C��7��l��J�%H�=x=�Cq��ޙu-k_pW}�J�,?s���s���ݼ�{���R9He��)7�]m��ݞs�q[�U��ތxou��8�-p����e�ڠ&t��d<Q�~w��܅��HB|g��8i	�RK䇮v�s1U��9���[�P~>m�P?�����aY�څv`�=��N�I륞�O�����m�R6��4���%nSIgFz�I�`�`��:�5">Iw���� ��:�#�-��	����:�τ�C���/oEKATj�~��x�buS�N5=�F�D�:�dU!���*E�1B�����Ҩ�w$�o���#�.�	i���i2�X�χ�T������^a���+K���MnӺ�n��M��w�[k�Z�0���1����C�/º9��\1-4���II�T#�+�љ�&Θ,=���ս�q߿�F�ZU9��ؠ�E!�~��a�����Zo
�,���.~��扨��6Q=���.�X��-i.J��w�+�!�V�Yh7��M�=�.�!�ɕ>�х�k#��&�MB"̷���я��V<�ʝs�9�U����kj����%*�-��MPs(y��]��'?��?�|��OZGS�őz44��X/���h��o�Q�Vڈ��\�;;�����ۨ֎�v��P1��� `� [��9�Q�c�c�������#���o�{n�*w�'ϳ4k��]����gO��������uR��?g�\7�Q�2 !'�N��ܚֹ���]��ܺe�$�k�� UN��U[�
�&E��-)H���Tn�CŅ_հ�E���H�6�@�Şb�`�ޒD2h�<`����/~�oB�� �;WvP��cI�@t[�R���������l��t"�T�E��ʟI5"�?^�$K���%K0��97�V��QG�.��r9�8��׭J@yp�a���M1��c{�w��i �h�qa�hL�����#�uc���1�/6�0��â')6�<���'bF ��v���s���7�-�~R��*u�C�R�!�s����s��5:����ջ����߹��G��0��(ȵpI��d1�/�v6P��{
�ޒ�(_N� F"����H�Jڂ����q�6UlcE�1%ڏk�p�2��	�½�m�}�INx'\I��̨SFbQe�$ �j�H��N�ظq�o?�s$:y����=�z��e����/��(b7pP�v6;a�V� ����8M��8�]��ֶ���JZ�B�^T��T ��{6#�Ѷ���ѭᘦ,◑�!�_��?�-^3�#�n���#��CHMuX�@�L\�cRN�5�M��5I��I��2i�������X��1u��ݲc}�K��h
���	@2��KV���`p]8�g���"���KPZ=C�+EЫ����(O�*ՀfЇ�c��o�	�38�!��;�b}� ��ə> ~�@�ܧD{�l35#X��0���_<���;���V��^Jrx�2reQ���k��7�p�[���5����W�7vҡ׬_�h��-���/���"���C��l��Vg�ae�o}K�w��vڐ�ЩPn�Wփ�/}�	!4z��5<~�=����A���"�����������,�_���峸�ܧ��Q3`��@E�>���x/<#m~�p����.|x��)���Oؑ�o�?���������^h���ʇx!��h��Ti��$WbS(�9�|��߫�t��o��X�j-�i[D���Ʉ\��p6��N/����ښج�AS�5��w
G��\�B�^﹈�r�* �Q$�Z#3Fu+$�ť-3=�a��X>"L�#��C�gP���~� 2>��wt��<'���yx��t�H�ѱ�m�m�v�#��Joy�7��mra�@�!��^ yr/��o�B\~����|ݩM%BE����:�3�#=�>]��ۛ���Ӱ���< �I<>�r���z�z�Зs�����	�'�n-�y�<)̛����	$(-����pM:2b���2vc��bNb�R���_�����o��ں�8�=����f���_x%|uϚ5˝peU=�]��U��AE��y_܉�KF��p�6��x�w��>(�k�aT�^�A�U|ރ���u���6��H����,��
K�(�u�x��餁�ڋ�X�J��J��r��C�!ߡ�_O���	mae�1V}����O^!.�Ӷ�T�)�[�DV��t����P<{��'�hC�M�P�>y�Ev��ﾯrW\q��1s����[��Ú��[�mU5:��8��r�UϮ];<���tw�;vn}Mm�2F�R�ֹ�J�E#+ڧ�~�F\��fw�A�ʌk����D����)ЎΥp��ꛡ��*t�n�b7C $\���� �͈V����f��"U��a�B��[�6ќ
�Д_�	1�'_iWxy W�����y�锇ϋl����w>! z	��(��6��ƞ�C��w��� ��@эrkVG�4|L���ǋۀ��ߣ��_(���{ 3��4l`)�z��>@����z҉v�rq��s��3 I�XF�)�,z�V,_:�������`j�TxY��c�#7w����6o<��d���h@��߰~�I���U���f���okb2
��0�;�dxC74���}���ǎo��(1����g?�'��C��	�����j��Y�z#�3��"�~�wLLi�l�X�6ګ���P8��0$������h׏��P~�tBk��=��c(�6�x7|H���9�x�
y�+�x��g�P�@��ޡ����Fe$Yz��s���Ez'���/:�K�^�k
��4 N�晪ں<���_������դ���ƍyC[[{�SҢ�9V]���:}��ҧ��.\�����-]���ߦ��v��14J���M���#�^��>�w���\+o�	�ߐ�k�> �D	��sэy)&<;�8Ȧ�_%����-�Y�ٚB)"5b�m``v!?��(8��N2�?(���" ѰbW
�hv�����wf4"��*߭a�o��?�j�3��&m���feo��� ��� ���K���	��v��$/�� �+�o;�dw�g/27��W<�>���j-3(޺�ĮԌ�r⤉9�<���ܴ}{W�x��r�]�m��9��L�tuA� l*͈c�
�u�;����l+dt�YD��^@�ݠ�����M��ڠ
Kk���yp��SR}�,�w̀�:ȏ"+i�;�� ���K��<C�����A�aU���G:�ҳ8�2U�D�	���n�o��)^����!~�P �U��B�֞v�;�	�r�W	����!� ���g(3}����������n�=���Y�����K��!Qv�7�|_��i��v�{3�?^���&%Aa^2�\p[�ZZ�;v�ٽ�}Is��Q�s�H��l��
������>�h�N�u:[PqӒ�$�X@y=�Uq�dƘ�%�Q�0儂��*�k��`q��D���aZGG��#�H ���g"2���sI����u�Z���H�g�a,`l
3Ċ«{����G����TЕ��E9��It/�ɢu֬Y-�@���S�eq�yi�o�)92�"L;����VL��1՟�_�#	��@���o�'芪��D� �pv�ڴ�|m�(���:�Xw�g�w{/��m�l~�Ε5�Ö��C3;�I�#]�H�x����2���ZV^*7�Qinz9�������M.�w�[6o�?4 8ؾ�3�<��pS�Ls�g�v�-RJGY�F�0�v7��~mr0���(_5�"��X���8j��`<3�*O�#��p�ƥ�hX���*��.p�+y� �H�lt��k@!�cpϏ�!m���(��=/Q�0Xi�<��Ƀ4ѫ��8e������w"u���׿����/����g�,�A	��ߡ/�o�N�P���wW�0(=��>��O��|<fc�B?�:�6�����I��)e���s_�Ǚ�g�5kֹ�|����dmg��i 0}���Y3۶�m}$Z�<���QnY��@-֟��wQ��ڪ���2�jV���\�b
\�(ӹ���k)UMp�z�{ӛ�h���Ԡ"4 �)P$�*�N�s�0��������i�Iƞok�H�8hh� �F)mu6�E/
Б�7�k
���xt,���N:��=��i����W�SWD\���AG��l�|�����g+�myNOz�I>�{��&I�{���3'�W�;���#�8�����i_��,}�~xR�A�&� Tږ2��b$��7;���*7m�;>�~�N�p�:����k�ҹ��/o���V14J�=Xm���Ƽ�ql?�|w�UW�~Mn�ܽ}�K_4}����t���1��@[��R����l�䶭��iT1����ǩ�y{�ho�~$R
FGұ�ꗬ2���;l�p��5��O��&O<�[�z�Q�5�AP+ާ����AB�t�8��À ��Q���:���Ω,��-F�w�а�$�ƥ�hd��} @��=y ����8<#�.�	W� �3EB�)�����y�T�Ѓu�ƹ6�_~���ww��wՕW�����HaG�.������|��2�#mP�bEhDl��U���ȍg����>*�=Q�iO>��jm.��p�u�}����B�F�mG?.^�ؔ��򖷺����j���;����W�=��P�G\ۨYA>/3�����ػM>��}�Z�^��~�7>Y�wQ���e������ܨ����\s�Q�{�ױ�y��w��4�c��g�8��FU# $�0�
-vD��������_����V�����PT��0x�@��i:�8af!:�(�ژ�����7H�,������	K�i�{�+&���?:�}�򯻷����_��Wv�4��^{�뮻ζ�i��jX ;���U?�rئb�P��WU|[C��c�%><��M�tc |:�q/u��S^ ˇ#S�;D��>@����裌��r��c�=���/P��V�[���|�?Z=�<^��w��xACQ�b\��\ݘ�/=�賟&�%�����G9.ױue[k[l�dӔ|��( �w�,�Ot��'����u���曭�?աMXg����;42�Y�CP�!:��E5q�|�t⡍���(
��ŉ<���.    IDAT%.�f�G����%Б� �b|A\���'�&�Xo �)_1��3<�Z�����zL�֬Ycu>���ݯ���hqp�s�,H���fР���o� �߁d[�A�E<��C/�6����L�e�.�����ϭdXM�1�#.�ǋ�D����3����=��#������K/�T���;�:���M����f̘ZЦ��� H@����g�Y�mx���;���y���l\�����5+����?���鞆3**�E�C�bR���}���w���E&	�M��j��y���f��F�q��׫$?4�P5�2��K#:�1��s��cu��z	p	������ACU��iO���r>��~�&O�*��lQD���ܪE�2ҭ1^V�D�X,�ʆR�FF���$�����~?+8:��lF�r�n�H�}*�:��a�%e9�$�<�� ����-\�-ƾp�76�\aWT4k/�m�%��LD{QOlߞ���Sqi/��x������\�][����fs�{���I��<���OD�5"$H�&O�T��K>1P�~��[��X֊����_���g��w�x�#���LM,&h4kD5�Q@�l�HTԨ�xB(��;5E��Qg��ޜ�s�w�w���T�$\{��M�qM�4�\�q?]k�V f�� j���#�'Lh���Z�l6��q�[�l-�>{/4C�O<>�tu�
��>����`ĵ:���L�6�\�M�6������%PM�mJ<�Q}�<� �Clk�|ł,���3%PV�V�
%fF"��hW�E���;��$?���ޡ��*N��{��xCפM]!R�3V����np��w�6�5�0H�������96�͛z�ڵ+���/˩׍�I��7i���p�5kW�|��m[#P_�Fcuε,}n@�i ��:���c�ns�Q�.�H,���J�ƯQ����6N$CEC1��kz�, ��x{G��� �iej����R���!��)�t�kש���S��� �Z�\��2`��z�Ϊ5f&" �C�K.�� �*��cI�Ԉ�59�(,�j�~®�&�ŀ�|�Ȱ�2��r�f�@)yT�F	��D���
�;@*vN�!��A͕$�`��q��<a��C�@�tY$C�#��6����GlL�XCm֌K\T[�',W�C��3r�F�-&L���k ��|O�s---���Ǘn؍��cO8���r�-�t(���sPǤ��8��JkQ'������� �dƵt�)��yh7Q�1Ѡ�5k�{�ey�,�'Z��qXV�#�b
%�D:Kj��%�R�S�]���̵�~a�:��r��J���+��j���n��vsO=�4��u˟]a�b���SO��ɛr�'�ʠ�J���nӛ��P07��lJss�V� ���
�ZIn �� p��ʀ���{�����a п��A/W,ā-�}ڇVD�mV.7D%���&�.�\���u�N���ļ�(`O�P(�т=c�@�ȗ��]�:���׃�����'�t��h��x:z��GVJ�U#���8�U���o:��LWϵ�._��~Z��8�"0m4m���\:�Dj�:ₕ3���l�dĚ&Ŷ0ʹ���$���h8:
j�t �y\���n�k=`�uWf�h�C\)�ػ(��1u��P���E����$�$�㘖0�=2T��Fٵ�I��5p�� 5�A@]&��`�g��α�خ��j{����[�� k � ��R��g����͂�z���\J�.����Y�ԋ��} +�I޴ruf�4����f��n�?����c�-�F\ڂ6�p�M�HV�vƫj�(��)t^K9D <I�����b-^��I�
.��y�-Ʊ�2%"DW�$ �`�k��!��Ih�چZ5.�����Phס�]�N$$HS�?jx:DJ[� 
�#�M��E�i�0�����Y�� �5���=�z�f���%��QD���1t�����D`�v0��pHhc��N�(-j�Y�1Px��X��Y7u�4��_�r�/���0��Ǝ������'?$K�I�݊O }�J~�5�-��5����@�FLh�l��%T��}Zp��}�8e�;��jfEzB��5��wҧM
��7�[j�0n�
{��~��6�_��K�ɿ�׶
돯Y��
]%	Ih�����y�鿘�J^�e���p��]j�Ff;������-��M�Ċ�)M�I��]�Ѣ�]6��Fי3�A�ӭ6�.��$^b�t��Ӡ�^	�`���(W���s�6�$�|�E(ZlZR���t ¢�GBj;�:
'�E���O��۸р#`B��� ���>q�JLG!�G�.5�p�#�p9Q^[�T�5Do��c�2XX? 0@�����= N�JE��0����g��ͱn�]���� ��/�-b�4mH{�1��o�f��d�(��k3"$^[l(y23M�>]�GcV��`�x�DM��K����.BQZ�\�(�\`�Fe���W.lٲ�$�R�������U3�l�u]}cT.jeRTZ�Z��h|,3�F��(T������RZ(�t��`�|&L��R���~���M���0=�e�K' ��h %+13�@u7]nu >N�i �CN?�t���-}(8~����<�V$��g���"��Pb_W��C�7�����كrM<�H��1 "6�o��)/�@�'�$ġ����� ���m���6Ȉ��A��[�Eۥ�W3'�����:��9N�1�͊��C���ؠR��I�5U�d,O��w<3n���כ�E^rׯ_���/)BY%��?�����mk�����\���k�xݢlw�ɢ��Ӷ�nk��a�ZnLݦ#.P�ǃ���c-T������f6Ow۶n����H�; ~Ş:m@i�((� ���\s�,�`��MA�+I3�Du�J �)Q�7J�g/�"�N�P���QZ �a_��݄qM���4��*�7ʁO�dJR�'�ڀ�A��ZL�2Q�4KH
���n����OSovq I�R_��.�jm�igX!�)j�3��0��8$���?���)������(�~�d�^���꡶�k�'�� �L̫�]/�R��J�T�֦�\B'B�$��=.���P��+�z�K�m�a̸�wvl+��O��{dk����������G�����/U���Lx��5���>h�W�K�To�^%��Ɓlv�<�j�.�%a�ĩP-�Z{ń:�[G�3�|���[Sʗ�s���/��\�Z�����h���AuZ..W�%]'d����fT�xA6g�~�m@�Դ
�:ƪ���_x��c�ug�u���<��%�?�$��{���c���QQ9ׁ�񌝼s�=�(ã�:�x}�>��Ύ�ݨ�҈׮]�.=�B��H�H�2�~JN�I�����%�a�A�U�1��)�CY3�|����O�W댬6��4 -�V�*����KZӈC�����O�j�:Y�¯�b�T�Wi]���:�oK�}<�7�5�*�>>ߨ��m��=���6+�+���r���m'�,�硕�χ�C�L;h�\�O�+���@�&��9V����+n��K�I�7Zn��`���c�ĢX�L)��EK���.����Tj��9�>����\����D�8քGb��3�ȵ��VJhƃB}YC]�ĐMn�n�ݶ�[���𗀊 8���y�Fu�>ޣx�4<.W�z�ᇭ<�8s�̱��,����B~�E��A�ZҜ�҂]+Td���f$�-7k��K�s���<:�����{�ԋ���Tߓh}��y�0�K�j���r�C�B�p#wYn�>QP�JKg��t�l\9V+�A~1R����v$uPO_n�]��A�#MK�������ܟJ[�=��)�
��w�t�#��Y`a�klH�/��/!/����&���*^{�wݛ��&��J��U0�2l ����;�t�ˇK�X ��qPK�  �C�����Pe�b@��98�%-���w<Pn�!Ϯ�7s�L���'#
e��9�`]����wG[:wĦ��Y,Ԓ%:hs� >��I�Q�yqsjr�y衍A��ǻ@���!�r�O s�����r���sҢ�ob݌-����X�G^�*,� h
�?|� 
�x�� 4���$M8(nN��=t)`# -�yo�	%��yy%~�|)�>�校�(Q(aӦ-�����'� �tI����*)Me��e@��������6Z��i?+Qf$�NKڗ)$"��w�+.���۟��%-ٖ���x;�m�s��Qn���/>!�%�}ƿt:�2c@�=�U7^W<8��AS=@%.�?,(	��|� ���Y�_�$] Gz��u&�!�ǳ���fj�s��@�.3T���hv@2q�%���@�I��!�!Mޡ���J���^�k�i��6R�F!��64��+
6 �u�@��o:�3@`�=PE�lPN(;ׄ�|���i���
p�C������ȼ�=*�lİ���,bаI��t�g�P$�:3^"RN!�Ʒ���N���/I#+"���X^P� hX$@Pz��H�C�uHC������"V���g��E^��ͥ�3��f�pq
� 0A��߀�Ai��F�u�*�;���b�� =q()�!�]���� ��&�O�
� ~�(6~���9Zw�"��-x�C����^��8����klG��B9;ޡ.��@�2V��^Ң����;#�Ϩw,�#q`�Q`QUTI� ⷝգM`3�>�N���`����߻Uk�s+�[54` -T�h�u�Mۼ	@n�YX�[�~;*����\!'~^�4X�p<��g�5!,P�@+�u������}�r�!n�=�k �8`�ts]+�p��Q%���pV�6i�^�-X��~�h_t@[ݩĎ����1*������`�s{�၏n۩(��FY+�o(���u���(p7�t�Xw̴P���Dx�B��� eo�%&]@�~�9���f�(��HCڥ��L���,ΦM�LJ��%�}X �֬^m�ed`Rn�3� �*�;�Ϟ�d��P�4����iaT��gkOt�����m�1$� &	�u��Z����2")�W�Φ�C�k!��֦�	�tmã=��
Y9���Gn,����{�<w���{�9;��qh+F�ZB��cD�v��}�_@��NgD���~kQֹ���H	y�d��j����;���[�l�kٸ� �gH�P�B�	G���ni���a \��k���$�KV��i��>�ܭ�-[�g�>*����%��$PK(��ν z
�̢�{H0��h����=��Z75���1��@(��G?�Qw�܅a�x�7Ņ�By1��;�-*��72;�Y��ʿ���u�]v�{X�6꿇�v�ʐ�2</���}֝w�y�e㝔t�}�)�g����neb��AO\��&��䟐q��wΰ��W��^'�C좶�D�@� > ���������Pn��vQd,�;�F�ަ�[���S����n��V-l[��>�Ԩ���M�ɂ�O2�3(�V���� ��<��Z8_җ:��w�˽��T$��,�Gy�X�F�N�6��m�̰!��O@�O �(�z��S�l*���_�~��IF�Hν�-/��Z�����X����"+�&��� �@Q�Q������Z���}��ƣ�����������S+�'d�7�|����0^�c� WI�Vj��e�Q�a#����tg�}��C<��O>���'-(qBJV�r2U��A��y��J !���X��Td)<E˺3�¨���Z}+JB�����c�] � ��7��K��Ve���;~�K�z�7����b���� �w���<*]f�@D4����5�c3Ė`�N>�++�ɀ���+\ˆ�n�[�w������T�N>���Ԅ{��%Y��gZ�SPo$.Vv�D���AU8�W��Zf���~��!�Q�Nb/�� �`TjK��'��ԓ �o�ov.�7(��-���7��	��	X���7c��in��*v*PR����S�-X�������T��z��bl�u\���3��ܺi�啒,��.W������vȓ�*�f�D��U�F$��Rht���Xr�ع5�N#���2�
���
� �5$>fVӧO����O�4��h��g�c�]G]���OD��%�#M('�� ��a0 Ρ.���0{�"��Sة<���߈zϘ1��J� 4���4y5]>�'��*���5����	�QG���{-HΈG55ː��+`z&�3`$ 5X$$ ��1�eцd���V����~B���S�.8�A'�4	l��f@��d��>��u�ʚ�ubs�u�6�c�9h��e0���E$�~Hh`oX� ?��=���Qg~�ڇ"�(:������i����r^��m8bDՏpaԁ�>�6�[�i�����t: T�5Ā6  ���o>�\9�����($�2*w���b��b�
wđ��H*��(�=���6��#�x�M��}���~��9�����_k[��v��@o ,���x���Pf��~
;���u�;��J�(���'�RuM}�������ʡ�?���x��m� l�`ј���1�@(�"���$`���|c'���*�'��B����jݺ{�<ȏ��/� ���s�.鍗�W�0?'�Ri]r�����	�,��gH[ZZ�y}�k
�>�t)y����y����/KUM��m��,�)���/�(`�Σ�rwvV�(�RbCl�� �e( ��%�;�),
��/��t�����X��J\��Ip�;���C�q�'V��=�N���/����(�9�Am�sf�u�������#�W"��_�t�׸f�(˖=���t�^R���aK&�V��Ϣ�:�3���6�uyf��5
���E�=v��˥74s� XP9~�0�
`��A�s3��L@��eҤj;7���i �@����s��c�I��֜��!�m}��GO�.%i�P/}�Q�#L�1l]{{���?~�>������a��Y�e ��S&ҁ-!P&� [FK+�	�X1q3�L�.�Q6yaDV�/u�6X��f����=z�N4�f �N4����Pp�s_.(��2 ���eQ���ü�։bZ�:h���3r�\%]���z�׼�xnxr �T~Pc|Pm��,qJ��:�Y�ʋ�"���&�-�T6xd��A'cK� Y���C��_�.���喊8��/�mR��SH?�t�Z\D��V�]�ϨdK�2M�ɲe)&����� jz�h�� 0P��ҷ���ϻ׽n�4��
hC�wP\dɲc�)؀{��'Lvλ�G�򁠴��K�kP0S �A:�T�=J�����Yљg���~�;�)'�b��%]�9(�^��w�*y�7����c��)�H����cN��w����-�@-`se2L�PPm��xx�š�o~�ݱr������&��n�M��0 )���CZhb�3F^� dM����W�#`'z��m��D{08�9�S��4i"�����/���c@���H��9����s:VDe����RJ3�����2V�]�ψ��K�MK��,&[�7@`�
���4x]��a? $ �j����S!��}�C2 h��y~`�S�'�m�3 ��<�YCy�� $�	�}�zSV*����a]/y�>	�G:@��;Pmf ����6sDc5X9�0��:�Npo�8 �U�j	��8�{6�Q��\�o��I2e!S�u�go_�͚���r�B��u�P <��q)���R�*H�����v���%����Lx�U�ͻ��|x7H�"�6�b/��_�FMM�ޑ>yF���w�.C����NU���l�ǔ��~ݳ'HM�h%���۫�����r�Hz�G���]?�Np���x����Aq�� �3(0ψ僢c��Vrf�ƍ7���GR�1�L�8��v�H    IDAT7&����2�y?܃�����M����rK�5�<8r�@|�!>� �0;q����r9�}J�z�2BGL�#�:uE"�f�yM���G���I@����6 ��68#�����s|�q���k�I=��qFώa�<�b�]꨸H�(���f��A�M��a-���,�`�`C�Kc� �8��8���e�.��������+g�x�n��[�'+w_^o���W�eg�W�Gz�����d�b1��
-�1 �J��D���()��f�
E�
��{(*T��p> ��/����_l�S�õ�܌��5���\4���т�5z!Pk�4R�((�ɡ��r'L���}��
#�:�����S��V=gqƌmP���ޑ&3��|����v"�Ê
�C�������R.7�dݣܲJ,˩���� ��e��6`� �z�g�����u����v�m�P_n�N��a֬Yn��*��N�6�އ�ت�K0��+�ѧ��W�����s���������t!�� ���Q,�?�Ye�����#�}��,ű��@}�:��� �M07åڈ	����/��L����{�]Jz0
� %�(.0A=s�����~�=����C�����9�'.�q�i��3|���gq�mc|�
s��g�T�0�
�xoX��UU㪙CM[M����}{����;קܜ2�bi��s*U���ŧ�d����R�	��i�1r��F%�[[ӹ�s"��4�8�� `�f���Y�@�=��.;}ޱ�b,
j��i������m� �
o�Q����o~�'Mo�aM���U�V�ռ�sd��*^�ޥ��L�ރ�6m�`,�\!�V��B���ꡛ���r�3��h&��{� ���Jp�K��qݸK(AY����d|�AE���H������v~����ͻ8MFz��I"h�Э^��s�a;�l�N �,6?���L�ì �vX|:�ޤ�D9ɏ2�`�r��x�y@M��C�>�F��O��Jԯ�%R�K92Z*5F����r�?��Rp7'$��PƅS5�  P@��*I?X����:=���E��ɍ�r��!��/��s�央���������Zy[z�j��轐'�JLF�-�>��������7q����ex��V-�\�6r�f@ןH!& r)��M���F)�kd�U,��IPP��/����a�sB0�7��?���N�c�9w��S�����:m��#���~^Rxf��'P߆����|�m��T�����A~�,|'�� )UyP{@��4Zo�p~D�lJq%�)��6�T$Y����m���.F�H��{��M�:g����7j����+iȾRȨ(S	 ���&��5�^owK]�v�}w;�]���i�C��y���FM:% �3j�E�
�<H<�J��$����}>�v	�kn�s(���9���=�k嵯�&�m�( M\Ր%ff�x�H<�L��u�bq[���I��W?�w�
�E��J��H<p��;(�Oj�}>��zx�׭[�+y6σL��X` ��	��7���N'ع�0i�'����^�V_� j�q?�P����q�v�[[��Ӊb��,rB��u��%֡"�L�~���6ʆ�I`ة$����x��'��?�+��`7ؒ�?�e;>�+��b����WG�J06P�z� AG�A�uO���Y�Qhv&���;�p�u�>�Ry_�e�&�enN)�Ydq�4@"^����G#����%����n;(=~�V H�X��
~���.���,��?�pw�G�3G���@X���}�{F�;��tD��')iB]aCB� ���oE��}���n��`�1�� z�D�U�7-���B\���s�Fp�_�$��E��~�'�C ��W|���zM�<���o�E���/��G����*9��=�AP�[����tn�5�Ɗ��F�mSm�i��-J��h	b1�9������Sx�.�f�x6U(i�ғ< ��N�1ʾc�}�<ŚT�pCg��0J�Mח�=��A0 x0���;��,��PrO����p-�Z$*nWW���y�<Ɔh���Ve�8�4��X
xl���q�Ȳ� "��T;���zXy���ܿ��H½�W�34�dJ�Hm!y�8�=�o���Q	�f�+E��82T��j��"
��=؁�@ƂL���5Y��g���K+vZ�� v�O����=�K�`����t���Eb<Qc:)X���X�{ޝM�I0�'"�D�W� �HL������Z�+Gj�_A��'©�F��#�gsz��� �`[B���=)br���b�|��^�nk�]�O�X�}u䳎���P�^�"H%��P�`^���l����@�Ȱ9��=�y���?���o���x�)>a����w�ml�� �� b&``J�)��.�=��{�w@�E��h�fMW�YY�4�t��	���C�<n|���!�KN@�(� ��7΂�="¨��S�dl�1!bE�5����٧"������ )"�^D|�z�:�æK��6�Z�;񤷺3���|N�n�4�d���o~�D�u0*���|b:�<�ʒ�)��+j����J�`	� 1�������à�:�rhu�7��B���0��ފ)�Q��_��Q�!��"�����������P3> �Xr� u|��_�>���X���E���_��TR�/_�V˘ �$�{��d%���x?Ҥ� �|��� ڂ������|���皼�;!@�0�`��w����vC���{SC8�ܥ�2�¨�@!33W���C3� 0P^
�*�>5 �x��ܹ.)����o��g�=c:�����g���ȇݏ~|��#uڪ?P��˔DR���PZ4�2b/����-�m�`z�a�߸�t�!*;�2]�B����}��K�}��p_>����+w1x 8u" l��:��1�KxR�)�}��C~�U�/UG�=���� ���xh�y��^�O"A�"/��� ���k�UW]���PMT[���<p�ZFܬY�L.���,^����	u�U�;q�̙c�O��)����ɓ����a�\F�N^,|��./�(X���{���~� .��R����b21aTR�͛'絃#��-Q����Ȝa�+np �E$�ڜE)��2��x\��)İ=:� �� �/��U��I��@ ��cG��QXʄ/p�_M^�Cz�U���=�'��)7i�<���\PtS�1��|�,��#(�JpK�[�+���K4� � 
((�� ��@�~�[�j`�3{�[��<;�:PȦqM:�}��6`�o&�ːg 6y�>��;z�\y�<-l��j�b�\�QV�y���_kG?i	�����=$@�E��wKd�3ْ�47�y|�ˀ�e -W@��X �"9�+T�@@	P8e���W���u������Z��w�o�p�Q턬o��#�6?)X� #��a 1{�7���<�<#j ���ǥ�W�
F�L�B��d4���%�F�>�T�V�6}�s��@���G#�#]Cq�I	v��� "�w4��2�����׿6�>�ܪ�N_������7$1��h6i�dY�<����y�C���E�Т8�o,yB���A���P77�4�5Y_^�u��R��V�j��0X(�^r��3�$F�#崄&m0R#'�Bpۙ���NG@9��w��QP���b\���\Š�nYڰ#�+m?΢D{�Z֭qW\q�m� ��%Y\'�~�NF����h@�� -�bO)��	f��k�� ��9���(�ǈx���l��MF�I�4JJ�r30@U��@�5�C�7�U��s���ߡ�sT2~
	w��(�RM����L�4��f�mSE @M0Ê �`�P��8�?����7�k|�X �����J ���%�m $o�-G(9��������{�x�bs��q�y��,���~�ӟ�Ye�]�~J,3ԝ5 y��Wyi�J�U��
�#:Hؐ�J�e���_G����Sj�����&H��\A�?� ��ȗqd��!�e��@�
?�;T����F͗�� �8q�Qq�p����G�1!c�$b<��y�)wU�9�dNI���7h��j7t�[��1�-�}{�vw����.���::P�4X��؏��zP9�W�A�_����x*�M��۴|^)�Īd��吐�aR�^��BJ�������}9���\9�e� 0��Q9��v��x�8�u�򖷘��I'��6h�/��3��#Pl�Ǖĕ���	Py����;�^z������w���E���Or�i刉�&M0��>8��#7�%6��а+�	&��E3p��7�{D ���EF]hv�ڏ�09��K�s$~X�q?���<<n��`SPl���(J?V�6Y-,�daw��xPu�3hx�4����M�[B|���̮_ߢA�^JW�R��"����o���9��Ӄ�׃��d��z���H����ϖ"^ڮ4�X���0*)���zmF�n�'P��n v"�y�t���dܘF����N�����Κ5��	�2(ؕ������%�Okq�H㩧�rϯi�"u��ڨ��.�E^�<��r�)�u�}��ݯp���o��Zm��R��+/� '��R�4pٝ�+��r]]>&Ǵ#&�Jpo�V�O�Q�K$������\Tږ�ڂemW���=x�*�'ݑ�ι����^�׆/�M��dQ�}L�@Vi j����Vz���㮷+�>t���S�~�uw��"�3�p�v�����m0��e�0�`]�'�v���)�LJ�Ȭ��J0Lf��o*�ŒD�N��L�$)ݪ��8�]Y�d�;۶��0���ޠ(UL�~��9�sg�)½��p�2˨�Ă�%���;+`��B��x���ũ�K��&����������"�=������xu%-L��ȏ`���Ǐo���	�M|t��|� ����@�=��<�m�l���D��g�zxgW��:pO���FS/r�L�\('d���et:�ۀ * A�l�e=,�@��K��K��J��q�������e�N##����7�!��k\���ɛ���뤴-[����֚4�<���Nw�]w�^#�9����{��$#c��z��d��l��tv�[�h3Z}�~zqG��]�-�-K�5RNE��VI�c$�u��j��t�$�G�O����nE�fW��Nω�'ϡ���PIuȦs:����KX��caZQ����[����T�k_����"TT�LZ��s�����]w�Ҩ9���
l��j1�f���t%���:[�º���ڀY	�f*���/�"ۚ�4�s������ۋ���Q�͛�����������w^d� Q��. ����η�==�A*�A0)|����NV\rl�?0��@��ء��ץj���Z9�!-Ψ���eu�:x���f�2��4F�6	����D����?��ΙG�����@�Im�)b�$�����c~�F���D��=<��>���_�!Kl�$ئ�Uq���!�30��p�d yH�g|X�A�y���{��ܩ�u��`(����	�	��
�>����<�#��Y޴�o"�M�6����m�c���G|h�6�[Le�]��#�x�nxpcY�P^�[rv-j��6�["I� Y~K�""�ۨ�vu͉L��>��}�1ڃR��Ϝƫǡݺ#��搠Lw���5�����;44��^���y9���{��,��ig2#�Tݫ�j��(� ������wާM��6��?�cF��]9���MD���0�LŢU#���$Sq��)=�*��g�J�#GDƐTTŉ�b��v�MV�K��(g�>۝��[�]�����.[�����i�2�S`{����C�PZtLP�x���M(e�v+�;�=���7i�4��B�o��;��xagV^{ݺu�!��a�抂�1N�	�(�d�	�����E?��6w�7ۂ�����9e#UB��oA[�|]*�j�N���xD6Ŧ���N<1a��[��u��~�S*�� `����d�P���^�	���<+��E�<���lP��:�v�W�8���;��Gf+��W�O\��u�Yn��yn����c�u��DVi��U�쫁ǢW�M�x�I"|8�P�/�%1�C�Ć����L��zW��fiE��m�\i��|�N
���(w��<E��Ɂ*0�7����$��_��W����A�9��j��vj7�{�ᇛ�5���܁j���<x؆g�%��'�x����Ysܷ��-W%������� �o��-���ƫ��=[�9�����,1Pq��D��P}ṙ��8o�������u�܈�RG���e%�<a�ڶ�� ��v05�3�s`>����k��.�:��G��jɣ���'�x�]{�5bn5pV���.�HMM���Y N���I�y��2��<��3,�s˴-��C��"6�*�|-n�<Xi���8��*�f�2@p���1�侴K�i�%C�t@N_��F�#(�R�-y�h��W �ȕ ���9�4��z$� <+���v4��O��S�)'�͜���u����`��G�Zs�5� ����<��'+��bTP"�a��ꫯv|�!�5ig����@e�kN
V���J��d%�ā'Ѫ"j�?�!pbH�Sn�x�3b[�v4J���^G+��+)Z��I}D�<����N-����4�ۛ��f��Y\�yƙ����=��f���}��Da�lX
���HW��J��Gu�Q^�5�9�2���v���)�O�	��W��v��6v��d�<�/��^�,�a�FL����hR��u N4�Hź�������V��W%%Q�,����kT�6 �Tn�2�Y8r~#@`��z�9�8�(�;�\���w�{F�0u�]c�V�7�1�q����x�������w�_~����Ns�Y⹱��w�}L�kì�A�ƍkl	�ܤ��C :��UZ߅cK��3D�1��r��n�=/?�����QJ���'WN�X�BE��y���C���hz�+;��$��5����-�P�u�ofc˜3�<˵i�v�Drx��EÕW~��a����Xޠ�A�Ix�e��o��s�=��ħN���XHH���{6�J��dU���p�qΖ��ճ[�bMT�WR��f��^�u�Bk���.l�?*���ԇ��_�JW�uؠcz�:C�q��w��3�">��;�x3F8��%^�Y�R�&H3n��FY7�"��gFJ���/h \�^��W�Q	��Γ�p�6c ���R���g?��QO�)3;�������L�H4VҰ��P�}�`C��ŋG�٣��'�ږf�̍ʻd��L��Udق���E@F/C=��%�@�˲�߼������|���w ��&
�����E�v�Ĺ�R��㠫MhsG�'�X�5ԍuw�u���W�po��7��u���Z�x�gW>o3I��(�m7�%�ں��xB�`�s��|��L���z�r���_�E�#5�4���-#�x2'&�ɘt�����a��w�n{��A�*����΁B� ��� '.l���z�灳}.�Bг1�]��l�d�yg{�(��� �/���'L�5O�΀op7�p���n�r̙;�]t�E��s�������u�v�$۲f�x�:�ր^��(#�0ȏ@���2����l�U�Tã���������Bp�ism6VG#%����~��%�\:<#�a���W�� V� ����>QO�shp0H�o٪���J���?c�N;�Ĕ���Ci�0����f\�����=���n�����`N6�o�$&}n}�����g\�FR��2��'aP�'n(๽��zl�ʈxH�ע�T,ǤӞ��)h,�\�Ī:"��Jp�ߝ�����RI6�t<����7T �lap A� |�J�X    IDAT �/}�E'*<�j��=)�W(:���\���fhx�4��[��^{.p˞~Z��:���%��K�R��W �.�T�^����?������(0�G�K]mM���V~"�=e'��C��pWWWe�\H�k0ީr$�.E�Z���0*��hM��3#=�m�<�έ:�`S���7�̀�ā�#��ꐤ��z�H�Հ�+^NԳ��^[��A�⮮ќ����	���wP}0-TEȉ�K�ɀι;�h
�� Z@�����m
E��n�f
U�����m�P>��ͯ8N2m�SbK��k��:��}��k�L�+j�s��;*���m�O(����JP��g Sw�uD��,9r��[l}�]W�t2����>W|r�d��i&������Q�-
���#}@K�Ȫ`�Ƣ��SNr���g�#߶�E:.���Rռ��K���X��6Uq Ȥ̼B �ؗ*�Q�蠺c\�)�e#K�W�����,�4�^��
   �^��%�Q]Se�.`d L���}r�v��߶�X�#�C?��9vO�����e��R[�C�D���G^�>��=���s>��&�����%`w�w)mY���� O�:ո��$�e�-Ly[��5�$�_T^�JD�P�H�":f���F|d�Q	�������6)^!���PR� �
`r��*,2m�Љ��Vt{�O����
d?D*�F�Y��@O�֘� j�}[�=K	�d��mh�f���w��5E�{{���~v�]�*�(=R��.��7���}�B��a}!㉼�#����#bxa\G%�{z&�Jݫ�>�{D�j�
*ᯁ���5K	8�?���G�O����x�ݴxh�1t�C�O��7*�����d��b]�.��꼤8�d�_����ϓ�b�5߹�=�j� ��X\�/WJ�-�0*�I�0",��"~�"wm�5�lQ�[�dA��m���(G;Ӊ�u���}�T�o��v(�R�P�p`9�~� *�(|�:E�a{[ �k��n��y�,�p�H�{����j�|挙���	b/Z��&���m؊���\}B�B��p���p�������D	x��x���|��|B�,!�Q=�aB�5�X��∣ޣpA�"=�MD�R�X!&�-E��|�H��NQ�:p	��[�n�֢��f���p|�BXW�~�Zyb�W�d�;O
O3f4�$�o���U^F`dA*��z˛�e��#�&Y����6�p� �f�� ����)/��<5�`--�k��-+�m�����@���h�>emK��bI#�n�b<k��#��\���Wv�0
�]WΥDBc�y���$l�- 0@���?��Sm ��T�������1�EC��矅$O��8�v�-[ni� ��/`��-�k�j**�Gy��K��a�`��=��?,���~�Iw�]w��+N:�t��ծ�u���M���zK�هن4�5�����Ŵ�#ENX@�DҒr$�b���ҕ]ݣ�Kd��G�X|ugGgj	�� ,�l DA�)�HV��
���>c��'���������vy>�� Jb:���(�?	�CI�?雯o�������ڵ����vBZB3˥_��ť��o��M��\x�%��/\�A5Fik!��a`�IT�Z�q�0X����$�B��T90��{�0B���NTNVf���>��PQe� P�+!HF  2n���=V�
h�����i�l�/7MM����x���S�E&�,,�5H�ee�9���PU!�Hl�ڵkm�g@b�U+WH��j�Y���!^��l0�����M�J�����BiC�	<��i��{<�'$��+�r<�!���t��0*�].W����
���`���H ����
O�>7� �W[#����Ǐ�`��p�;��8��)�`Q3V������ g�˳ �h����cB7E����N�'�|ܽ�q�ۦ�(OR�,o`�pȃyT�AI��N �a��@ⷼ^u�;�P^�dI����6��=ɷQD�I�SH=T:�Ѐ� � �~�1`Y����D���^w��6e�[�f�tLnv���&��B���vx��`@v��C8w� ������9*��:���w����̠�XD���y��?ވ��	�)+�����������%�Ή
Ҙ�೬�93����	��r밺��i�bNC���R��xa|{���7c�$���Iz��9�Z\WG����ϚYF	_��W�;O}�9��?�,�$B���\^��;�z�������C�VEnDO��I>>k��֥H�X�-���5JLR�Vq���W)�qQ�I	�A�`����w3�f6"����LjG*��D^*�LJ��u�{ڴ���֧�W�Q(t�;���HI��~��3�k'ˁ�M7�d�ϐK��+_��[�j�m�j�'�S���抁S�8<�c���X�����Ͽ�����c�<�#��VF�LZܣ��7l����!����q�/.��u�Yc������5aԁ;��Z(�38�7F�5⇽~���NlE�:�~��6/j�V �wJ[�Ȥ��Dj�6�� ؂��OMZ�nI�PxB�;��ʎ)]�]��>V'������Z�v�`�}� x���� c� �0H������d�5�M�T���rz�܈�Ĉ�H �K]L[0����1��oѱ��eB��O�^� 8��$ ����d�	���X�[�#�wJ:��GG<�@�B�|�_�e�=���҇gl���I�SO-s��|�r�����WK|�x(JawI��@�\ ^�8~0���&�^��������.��bm�0�G�lD�V��;"P���,��5]��9\tq^,Q54�B����0��zV�<Z_�M��X�3�M&-9�E�/}�2R@>i�d�+��pw�_0�w�j�������;L�5�HR���R�ɓ��N'�9��a��PZ_�hZ�����˟��[����U� = �+�D���*hs>���W3e��R_]}�vF����Ė/_.n�(��v*tDr+n��	���v�g����S�W�F'�Ǝ�wR����y�m)��,������2�3�=��$b59���O/�0<<_u�{z��ģԛ�r��Xr�d2�)[� �$����P�ԒE\WW�{����<q�D㛡� �<�Pf�#�8��}�<� P������X�2��T��n�͞1h(#�D�-�}��J���#Ik��Kdzr�����R>Z[;��;[մ������n�xi�-X�t!� �S����K�5p���/��%��д�iӦUikmm���j���:M��������;���H}~���'F��I��hYs}1��b��Fr��&[j΢�1�.h�!Y(E�3��HT��ڷ%J�h��ݚ�d��մ;�ر}��Ha�<`6�S����렣�u�ف���G:�mj'�@��g �k�q�s�"Ӡ�o �I( �Xe�����^:"8�� .��	����4Pa,�E9�/$ZdJc�|�0��ߋ�x�K���.�ރ-	&�s.����	0/XZ�+�����-ֵ�u,�0cƪ��{L�Z*56��*�&L㸆��]9�ɕF�b,���)�E92k�>:�-�(F��h)Z,um��j!6_��do)2�M工]��N������L��4���6�reK����Q��K��������6�4�Iɪ�"��I�a�H�8�*)X.�uu�|Ok�:^��R�ڀ蕓�Bv SǙ.�BNjrZ�E�E�S�G2����ܪζ���J�\���6։���H����	�C����/O 0 pf(F�� ����I��28|��OVD�H. ,:( 0�R���-Gq��2Q��T}܄q2W�Ii%���Y�:yse���%�	�b�.y00��.�s��M�ԋ:�qݫiH�^�d�ɾ��f�ŞX"9X��z'�tQ���II��"A1���"b�
b��IR��~����b��:]9����<����3��L��*_̯�<����n���C��j�ͷ�?�����/�u���x������T$�O_w�Q�xdL��;�l\?`�%۵V:�¢���v��&W}���޾�v��<�eiF([H൰�&�^��b�!�l?ƻ6`֬��^���
c%,@a�����H�:Ǜ�������5#�[����*�:�ԩS�NUQ<�2���f�8@=tY�G�ճ{6�@2X�fx!�3&K��1 ��wٝ�^9�L,ɨ,Ϙ��y���`Io��r�<��\���j0�i�l%�A�,��d�Rn�����~�G�׽������%=V��l�rC��(e����?x0s�ո���W2����5�!������O��W�n�<�Kc^�W��ԳJ�����ҧ�N���{�{gwe}ue���{�ޓ�޹ra�����k�o��{���ǟ���o{�;~$�~L�����>�03������W�f�F^�v��3�7�����Np0�D�Yx�T�B4��R���	�m�S�N�2�A�uu c�g:S�;�B!�⊩�ػKj/m�݃��	�k�W����a ɿ�7�F6�����S�xO�L\�O׶��]_����.K���ͧ��{�~������o��L��#a��sr���A��{��*����Gԉ���Gg�����EX L�YyF,�����ԭr�����l|�<��U�C��O��4rG|7��Çv33|aucm�����pbym�On���>�zv����?x��Gn��ޓ�W&������<���x+S�^�g~���W>g�Z�gs������qi����s)z7�{�H�Ă�xn6�n�,�c(̍��`!d�"���U�3��/��o��L�
D��`ZK�)&3����~��"!w�E���΍	�$���������ۓF������w��\V=��X]XW�g=�Y�O��O���7}�7��Q�q�1L���!�<]�gTou.���ׯ�i���3�z�6�h1�����i�>����s�v���<G�-�w��jYc�{n]4�����3S�ֶ7ߟ�y��������Cǟ��C�����2���DV��Hq�K�No}Fv�y���Sw�̎��DR/L7�/��D�/&��:�b6�~�U+�a����ǃ��Pq���O�;�R��.�e��N�C��75૿���Lw<'��*���E��QgP��7|�7����������g6�	P�g�:D]�jF��Hy�t�������������u��G�o��p���aR��]���7u#:r��5|���:�bp�ŬE�z������mu��0F�)G\|M�e51�g��m����3���o[�3/�랻���ͷg�^�s=>��=�O����������/���z��>|`!��r����;T� I��w��t)��#&��Or!;H��Lg���dt�٬��q8B�D�`Vя�2IKj#:�C0&�lW�"U�T�N��O[�BMZ��ݭ`g�+}7n�t_�z��{�Sy��]�Ƥ�Ν���7���_[�8R��US�����V�!�j�`"���o��᫾�k
�����L�	��7�����8Ĝ����gŽ�/���d��w;a����dZR��x��eSc����kX>������=��c,��e-�L< �����SK�/�˶O��?~��#7���>�߹}��F:�� �@����0w�7�n�����寞���ԕ�g����9�ըU��K�d��[���b<�q7��}�6E�q�+B�Q]�i��t�ē��(�܉�Ӌ�P%�:��]Ҏ��n��<Iu���OD������|�v[�k�s��w4.��g�X�q_6������B4㊇Y<;Ռ�ˑ#7�����,�J�.���շHkV�ƭ����+����о�M�p��O޹��ңw`R'��r��ā���3^��hc�ӧ��?���x���?�1��dm���ý�ؿ�����{M�bn��N��~ڥ3g��?w!���# �6KZ"*�
�ƶ���9�T�B��;K���A>� �"C@�w^��S���b�j��Dhy�fR��H��oٮ�7$GD���,��Q��vT&:��$�W��e�{ߜu��$Tҧ�t/2J�q��+��j�H���F�ǳ�ál�Y�@}T�������c�>�|1qMjh�)w%�U�:13���w�޳z��X�g#S6��L�*�[�7��� �w��מ��~�OT�Ld��"����h��d3�&��˱)b�Q��r|]R畩;����/�����S���O�m�|��<<�������0|��ӟ~iz���o�\������?�cͨ@G$yf-�q�K�Z��C�|�h�?�ư���/)�FD��|$�W����V��C��nx�w�S*�0��`�%_�(ґ�&W��]�ӧ��x ��ߪ�ģ���W~�`��>��������8����2��˦��F-�����|���k��kU���\0�9��J"+�[�n'�QSTM����u��W�2��O����4�������)=]�[�}��* 
p�^ރwf��OV��fvh�!�ď}qgys�O�f���>r��ҍ|8HO��c&�����|��.�^�ҍ��ϟ�\�5{I�ؿc+��h� ��JAߐY�a6��pQ��Z��$�3d��^$��3�l$'d��J��T�+m{���f:3�i��]HL�Uy����^>�'RK�����NĢ=��|6�l�c+G��XC~$֍/��/�e���%/��bd̪�$���U񅬆��c
| 5����V�=)WL�Fz��ɜ�v2:h, {&�1f�\Iaeß���uBS��ta�\��q�L��oA�ɿޥ�9ݪ��$���v�2Ѻ늩{��U����҇u��/-uI��u��v!+��8p��FއƛQ�&Z��X�,������}��Ɇ��0�ߖ���r��G�6�"�E>���W<e���?�Z9��O�8�"ڎ�{
Ѻsā���QK� ���B :e�뾈�u���� <��ż�!����K����K��Y@���C�I�Kc���7��~����S�F�	$=��bz'���!P�Yx@/�c�����L�R�^����^�����ۅ����۠W���V�^�՞�U�JH���R�s�+ߙ��{x��-��<]��&$���|U��$Iǳ�z�Y�2F*���#�mrh~~vcb~�������ڔ�UE~������b~ߞ��W~����^[�x㩓��`�XWX�T	����V���vk*��׆ i��k��0o���֦�+$�N�����e�\za!oļ�������W�z�^�`
֒^7k%�C�>��R!��7d�8Y_X4�k�8����eԱSgN� �0�`
S�/=7�I��߈��p滼{��꩗LГ���;�*�w~p-��4*��+8���iq����^~%�o�kKs�z^&�X�b�Z?t뭟~�����>z�����w�N�ϋ��|��֗ޱt`�;Ο~��# r �Iӆ0�O5
y�!�*�\�#H,�.�p���+�t�.�K��8�}��l.�Yߣ�\!T�����o�3�]��|]����l��ggx�6�w!���<Lа�aYN�n)��m̷���K7M:�.�TnjU��G�H<�G���ޘ�6^ة��V�����D��+������*�phR�������N���Rz�v[���S�J�P���/�6?{h�����QM�|̘��g<�kN����;!�� j@7�QsU,̑z�@��~D�o��W$J���Wi�����Y���&/i��iDH^tu����C^D�W��ؤ�P��nԈ�&eC���1Q�9�}+u�٪�F�b��=��R�t�+9�4J��w��#7d�Υ��rąem�\T���.:�1&{cd�jvz�'0Ի��`���װG�
�����z�c�!���T&5�Z�v����aΡ���A��[��QgzV��qYp�!/�S�
F9$��_$/g�onj�ݙ�[��6~>ƈQ��œ��1��g�����y蹵}A��Pk���P�{�p��|�
���uDt��Q���
����M�;�i Z�(    IDAT�A���z��Ȇ�$����J|���r��<��~�JJ���w��T����ʵ"G�����5n�6ÉI�:�ݷ���:^֕G�Q�]�����R���|�����/�o���U�����p��{5sv:��a��Io�y���v�1�hf\�^��鹩����55�I�'�$�>&�}��Ϻs��cߟ���ni�R�9��u��{e�G��8.i�M��ّ[�tŝq��i���l+MbW���k��"�����Q��J�Ew���mq\%F4qH��0��6�D|R��b�����+8��//s������e1_``*4Ѕ��8T��Wӝ��$t<�����_%���dV�[ƣk���ge�O�j\���GȢ�<-��~י|���~2UT���V�-d���&p�A\i�+[����ixe?5�rg{cnwfϹac���6e��D�����G�.^~S/�q~�;��f%{�	T�.	 ����p��&qB@i;"E���tfw�w?�;�����g/��?]�5¶�:L�)�Y+�����K��tkR��NiH�Z�������pI���]:eˣױ�������4B7��o���o���=2K��ǵa/��_�>�wX�������Ckߥ'0�(��峇8A�<�t-�>_��>z���{����?�l��E7�U7�RKn�F� �WƳ�{'N}+a�/[%1is�W������S�x^9N<�z���x�ίK�e�.ť�^7N�ҜU��!�t/I��Ҁ�RU�Ґ���t�M3��}��W�u��O���)#ϥς�b��!ӣ|{�������M`(sq��.��ΕOz��oD7������������|T�2UL�|`wSz�C��D��HeB�D����j�=��"�dƲ��#�%W�������/6V_nj]�p�h<K�5D^y'����<��Gs߉wm^��o����w��w�(N'��n����0��4=�o���u���¤������?~�������p~�`l�Wur�)ӕO����^�t��`�^���^�w�o��;�V'sgcF�{��\Z�A]����=C93;w����ot���uC�EܦZt�_AT��`�IZ-4X�v="��b녺e�~ @>���y׃wtY��`!]�|U�k'-�밺�!��i����Ο^��ʾx`xA��_@�_+�ʧ��I�OX����
BX������y9�<��奣��������o~�!q�K���в;����g�l)+���`+��J�ȧD�6s���~ol!n�t���Jp���粠U�������&�o@���7�ẙ;@lB�[ٚ`:�P ���u�"W(/n�<C|W�C>���G._z:��8�*XZYWผ�In��iy��c�������~�
~k
�Tp���T���_O���
�t؞(�eX�m��v��zW̗:=02�:�ۜ������I��No�@>�D+�.Nm�f��I���J}�1^�N\�����a}{����ŻS�Gt�^��j�[��|Tq�_˲�n8��xTP�F����Ō�B]�.V
�#f��t���g�]�B����ECZ�m���&I+�|��fr/���t�K�$��;���D�~$E�)kE���X�Ȋ��F ��2���K�$��a����^a�n�zW)1�7����a*o���O�ޣeyU�'��U�x����l�ٟ���m��2�e[�c'ZG~�3��~�r�ک�d�R[a0���][w
[�5llm!-�OV�e�#u�"�ɐ�s�{�O�$�u��qM�^��	]���Y����[m���3�8rլ#\����R��!@Iki�$�������/smp4�,Ď��oq��v�{�2�n���'ʣ�8�(#�5䤪t�6�+y���z��(���0����c#f�7y����i�{a�\��Bُd����'}�'�5�B$�ox���t�-�Ui�~{(��])[�w
���#���Rv���+��
�v����K��ܸ�a8������2���yt��<�,�+�?ȮB\1�HH�BР�������X�;QZ-���1+n>U�ѻ˙]s#N+3�b��E�� ��	-�����S����*n"y�ǳ��ӞG�I:娑 ������>W\>���c�	���*��Cj7f��
��Ԅ���ٟ7<�YώE&[��-��ٟ�%�4�C��U����?��/�Ҕ35|K\~9����邋N-�_�|HyW��\b���'S�痟��/�;��=����u���{� �<Q��^AxG���W$w#gϧ"��H�C/�?c"i�u���L�zz�����ǻg�����Ov��Fx�l*��\O�g��`e�k�ӌ��^�h��HZ�z�)�;��ӑI�<�7&=�0����o�NX_U4r8,;���re|����Oy�𲗼�xA>�eU!��tT_&o��{�bh�ǭ����w�v��<=w�0\"���$x���ލ������ B���s�v��Y��X�߉Ț&�tˍ�*���@�˱�D-;������t����F����� �'`R3��-Sl-JqE�*�Z�^�	2'R�PD�UR�Ce�Q�'{w1F�[�3�[g"׺/"��K�[A�).���u�[?�{�<�7��I�G��+��`+�_;�/��78��-~�"e[)c�n�")W�B��tɊ(�O>�;}����9ab-�3o�M����l5��j�疲�KV-e3���f�c�����d��ȅ=sSi�ᡝll������le]ힽ{v7&��H�'���q�φ [(�iE�0g&�;1��A����K6Y>ݭ��� ���p[��(����G��2���B���9'q�tյ��*�����yYjP)^��W���z�Ԧ���=���ɫ�W�8N�(]�Mcz����p���匿c�06�%��Y>�/��R��v����<o�b5��:���UY>��ʋ鱗+�1�U�����O(�I0+Z�VC`���?���w�}�����~�44�Hh��� 9N���K�-Z`�Q���C��U�{��W�5^N/�U=�8��"��s���|#���Kc���c7.�\�ɵ���/M����h�ַ�0���n�_�ɷ4��HW�IFI�]kWhЭR�5(X9`Q	U_i����#yE�,���(�3�����7����YN�83<���*Y�iVa7e�����q��;�=}�r/n�ά��	:�$�9����VM秪�F'T�2��y��?�j�ܽs��/�Zd�W�(� DjAL��;"X�ᣡ8�	�[�b��#0I�Gtj�@��������h%y	wm��������-��w��{��(mO��G�}�KO��Elq�o��iz���޳{ﮪ�(^�#RB��2{��3ّĘ�ۦ1�{3ҙ
��=V^����7�B����+��A�͑���޷��C����A�dJ��S�;���z����<t�(��v�&����uI�ai����LC�4��q�w��_u��qF FB�[ġs6_UJ|�5$f���(u]��nZWN	��o�����<�7I��z~y7�OF�p�W\���@Z6�|�1].�*1�/߄V7���Q.�6�V�eN�kJ��N__|m�h�ԓl��M�,���T�����zD*�z��g���������uE+��.���C4 [6鞼�?���[�!��2f�xs�������`0桊�-���8F��Ȏ�Y�=�?\}�	����
Na����r�� �E��Pg��w��7D��->?�&���ɧ�����z�^;�H�N��siE�_;�^uj�V��}1��}�?�P��5p����\�~8�zZq�{?y�|����ԇ����gy�����?���W�Doy4�vOj�te���ј�ѫ�Ԫ�ұ�����]��d9{S�{����I|���|�<.� ��[٣7E��Å���_���t��U��b^LӃ�l���k#��smU���z�'U��J�w��ܒ_&�Uy����d�sT���֍w$���t�t��x��2���7��Ǔ֯O�hT�e����W��wqFگ"]�/8���Xޏ�<��n}�Ϋ�/t����H$��$梃S;��7�r�����=ç��u��z��p�Y+�y�_���Ut���7?R;���B?�<����x��Zp��=�,i��!a"[q�15�5mj":C�$ ?a�Ȭ��I�^�2lڢ�v�t3]$� �*䏈�s��ǉ�5Jk�pa�+�������?ګ�������0~�߹��������޵?K/�x�=���ӈK��W^��}�Ucz�^�g��w�{�����y���w��S[���{�N�<�#��;L�����d��w�o+5&��7�0��>�t���I�Vf/ϵ���a�����'�V��������LF��%��޾�{��+i=Lv���H���uN+s(@�y��ԯ���AcBH�Ii������xR1��+�Qِ��	ʰ� N@�N�'Mu��ֶ;"/K�Ә�f�6���Z���	����R�*[�|���;q��
�U(�Ӌ+�n�F5������|*⺧�A �ŗǇx��b�.��=XG�;�f�>�t����/�����o��on�	;�]#�-��l��W>�S��G��*{��h�����@V'͆�eUJ��V^���~���[��o�R��~fI�5�-r����u1�����`۾�� �s��*P���>�|V�v�g��p��ϛrE(��z���ؒK��8�����`k3�b�c����d���Gq�OB�LCh�{:�́���K��^���myW�����\]>Bj���z��Cބ���j��J?V����B�{�O�1���W:��!.�VY�)sq�ۛ�����~�R�߯z��>�/����}�p�����~�6���~ș8Q˶��%�jS3�'��Өغ�2<���,ip�Sӳ�Lޝ�3���Ԥ�n����m�H2"r.�B��m+8r�8�I���"�c����b�D�-�c �{���þKmr!��!H�=G��<�G'�&����-�M>�#��廸���I�&)�=y������ڽ�͓�����j�����_�Yp��P�	L Ʋ����Vޣ��>�t�}�~��|\͕�ا�έ�ɉ8�|�K_:|Ƨ~��-����=<��o�v��_���ĩ�ɣ�䟊��9`�p8=��,0]�eñ���{���OfӚ��L�'
���'�>���3�eH��T�%t�}/���uƤN ���J*cdӿ����B���!��$4�F-�1��oN�9yY�W��?O�D�
�+X{�L�b&�UNoT�`y����������)�P�?J�����.�����O��Qo&8�@�D#_���UP}m:<}H�K��;ʂWe��.������k������A��S�����=ï��~��>�6�ptq�[�e'��ճӣ�������&��ԫ�0 K�o����(���h�_��.�^^>2�8s�� ���( �����}��	ө�|�y�
\Y^�s?��>�ޓb9@(V���oz��7�u��}�~���=o�ɟ��:�#,.�+��ʸ6�r��v�Gjh�z՗�hl����;�����lͭ����֒��	��E䗷)��1��Y_Á)��P��z�����^��ڜ�.��?tl����:#k|o~���[��IɰC�i�(<ZA���v&z�s����$2&FGA#��3��չ����z��/��jHg�س1���_�_;�c7
�������{���a*k)S䰖<���`l��q�F%�]㣚���S6b���'h��N��ر#�w?�  H�!oT��Ґ��g�7�rg݀mo����l~%vR�:G�����[*	؀�U�9s�B��;|�w|{�Nk���?�#����	���ј���{�a��ī�+��+r<�E`�����J��^�A>���J���l�:��-��]��L��ٟ��÷��簊?�?0��/����_���b����3_��_>�������2%��0�������3)-����*}7pe�y�q(=���՜t�/����������-�Z"~���_��_���0Ҝ*��8T�ip5H��aS�{ev!���q!0������1���ܟ(\��a�;)�rP8`��X@b{�:�L-���Ib._��_��E��d$�{2�0x���}��8>�s��q�)i��HC�k%�r�,�G��޵o޷oms����^���d�_�_P�Ol�Ԇ�V�W�o�=��՗���>)�`r�]���O��=�)���\��;���%a�����;���m��.���ۯ��a����ׇ���/̱#�~�~��%Y��K��8T�B}�O�upO
��Fk�|3=�י��gsϥXC��l���a��g�<8�����m��c1���b5Qi�/���S�����-��nY�S驯�b_�3�ʋ�ȝܰ���G>�3�m.޼���� Pq'�K+@���y>[��ǜǬ�mo{[I�8����˾,��;r��㱶L�|�wf�ǿ�3dXItϘ���.�3�z]A`�
9�k���B���g��q��|���~�T$;��E9�:�����g���\}���r�9�I�w��g�D�x��v��������C�E �x�;�#Y��ַ�%R}e������P��?"�_���}o�+Fcʿ�Q����v~A��u_-�����w���Y�n�������E�F��,g�:9�J�O<�p��7���Anػ�+���iП}cL �&��}�}oM�ϼz���7g	[�2"����?�����?�;<���°�BL����W�{@�Kna�U�+�>����4����>�6��ew�ts�4�o��?���I�?���5$�+~���3�п����YHW#�82�V�Y��&Tp ����XjFk�d=�Cf:i���Dv��xu�ո�y���Y7�gk�����#Q��ﾲ˷�H��h���3U�m��#=���O�VNb6��ȍ�2	b"d5�|=�g� ��I\sX�c9~��>0��������^�ۤ��^�d\�V�)����k���M{΁����Hە���4��Q/Wt��������<�T�O��ό��[�\j�C�X;������7���R��TK�Z���.��M�W�I #^�f!��ɩf`m� �r�>M-�IO,%�'�yjT���_��+�W����K0��6Z��A%��ظ��a�GI�d\H��*��_(�6�7���&6���w����_ĕ��ѸH��Bڨ����׿\5��J��,?ݾ2�{�Ǫ�>}�'>88�@5p�^V�zW������o=����ܻ
tp���A^��J6ݜK����|G�Ͼ��/��M�U��n��v��ʍ��F�ꃦ�VWe;5�۾�j=�|������f)o:rc�{Q���~���9��Ï�~�A�B��W���~���6r��Ɋ�$�.�I"=�������3��;�DǛ/(2:@4���>$Q2�,W��BN��� 9J<ibU�D>���v"Q>4<�O�@�͒=/Ӿ�rP�#a4�=�z�S���aLi���eԔ.�FnJ\�����[܂��`^�o�G���nd��/����_4���Q�W^Ș1��).�	�|V�c�gd+|@@���o��OPʋn]jNf�o�*������/���w��� ���k}��~�Wf&pf��_~Mj��z�R���
�wW�m�{Ե������
���c�Y>�s>o�_��Ұ��ON��3ܐ&��<���{�뻇;��$q^����4|��}M�ٟ���͎\�p���1� W�Oj�?��)\�sOM�9���r:�v��ԃ�x �k�u1���R�[�,q�}(=7 u��W��v�l�a��� KE&#-x���^R2���l�^��/zQ��㮝��Ï>�ٯ����1��e/)"p��������%��}5�Q��'C��i���=WL��c�����%1������J{��r��w���QJ�!����=�V��_��Q���    IDAT��n����+τE������ַ�e��O���<��#�Z�VQV?��O{Z��Ǉ��h���=�%��ww�R�w�F��O�Hh����j��v&����e�K�6��~��_��_�l��^=V�;I���oƔ/]�bXLj���P4��zFǏ4&ox$l���o�Lͦ��i��̮K-�0��r72?��|��g�����)M��*�Uӯ���Ga9�2{���
�Dc#G��w�n�P�|K0�I�\�<z�C�4"HZX̠o���n�0��$��BL�4%+����_ؽ~y�K���I&?g]�G�!y#�������� ,@ӿ�Ù�n�����Տ�*����dS�R�)��kȮ�<x
]��wy@X����g�}�;��[�7�H�����|ӑ�[n����� ��F�������B���58e���3�4h�0Q`h�a%0�&ϟ�@���kH��	�ӳ����������wxg�"t���i9é�xb.6�c����o	i�S㔎O`�(���[�ի,_��y���z8��1������ǎ�i��/.�wI���%v	٪� �Zu���c\���m���5*�;f�����
�Or�߈�@Lg��wI1�wo�C�u�a�~_0���gc�f]�?���CA��p!'<��廢,?>�$���<Z�1�ܫ�?���V��	�������W?�_�x���w�u4=ȥa#B���MpX�63�6i~����п�|!��j�,K��6�z�k��_�Aazk�&�^�������� �ıJ/F׆K�DW�xG��l�܋#(��zF��3�$5pV��|{��\s��ݙ�����(�!�I%�
��ݥ��{3=�ƞIdȃ�MDZ����$����gϓ`��ݩ0�ެ��Z�r�ﻟ��&r �#���LcVVkdm��۠���t�X!�8��m����{-�*ǩ��6b����[���x�x�.~T�b:����H�{ۼ=ߚ�.i6�A43�:a���������O��텃��c�|��7Ǔ���G�j��kJ�+�yO5�o�U���i��L�����>b��9ٍg�k^�K�'dy�������H5(0��� [����(匟sΧa4o��l����IŏB�Uc��O0eNN��(X��ӱ�go�ƶ5���듄���|�ȯ��dN#LcQ`�ӽ�]G�g��C�F���I �2C!�OB�=�:9$� ݴ�]��U{�a�K��A5/�2��_���3�,^�^Z$�j1e��^8�'V��4����P0X����\��-�{���v�v�mW'Gj8���=�B��oP�"(�4�*�Ӆ�Ue��Ry+��wo4�3k��yz^m1Yv�������a��/��r��+�\]<w��P����ϖ�O>�\'�6�ԊW8����N���A819��ẘ���ޭ�L~��v$�AGH� ��R�0F�f�1k��vk�Al���a�و`�ࣙ0�v�M��t����2X���ЧcT^#r�F��b�eOhAtG-���J3B2����Ԣ��at'�Y�D�Y>;�n�r���j6���9R�zT��p1ug;/�>_�m�U���I���xR��Y'�k�Pꍾ�#��<�0k<�K7��TX�@���icN��վ�[Z��<&g�ங �0<p5�쵿�_+�_~�_�A��	g�c������έ<=�\��g�Q*'|�� ~��Ō�0 �M��Z���a��y����#�6��O�����D�k�P�0ĐĐ��v�&���d�1�JBZ뮚����#�H)��FD�+���a�^�RMO�>dq�ԨEy����Y뗆���̬�����c�vG]��O�!Y��zzj��"����A��N��/�y�H�yO��t*�qL(a�����x���𑴘�`� ��#�yYL�Ӡ�.x�Ȯ�c���0��?u2L�E������ޙ�	������	�ݎ/Я��o��M���]Ϥ�r��0�Rz@y1���2�3����'�����mI��4PyD�f�Y��[�0Uë�\/s�����V��R �}T�=qi���:~�x!q&-�ַ�đL�$�_J�O��v�g�T��q�Xf�G�ϓ��j0�/	����g�K��0�l'`���{C�W�1�&�WVNֽ�9�Ue*�85&�4ճ$�Z�Rm�qb�|���V�_Q	��`���J����d���f7L ~����}����`�)��1��W�8a�8aϬn�\��ܘټA5�0#��;����lcv�C�P�E]�7e}$�F����z�a �F��H5>��b�:w�lᔰ��	�C�r͘�"��N���p���Kq�:Xyj �"�`�Z0��PL¢g����e�F$�n.̡�ui� h��fU���~v�������r����R'}h���r���v+]�pVSS�1WL99�f����AV@��L�t ���c<�Y\j��z��c��`�����5k
�|k8�BzoԞ��BL�9�0;��j��Y��1&k�ڪ���Az��O;))��.D�.=8���2��`����$(ݐ	��;��&{ab�$�3��BL��w����1IO�b\j���ķd'�����N�lG�۹��!�.�A��Ԑ�2�_T8�j1@��աzb[Dx9
�}SW?,����2w�ڞb�Sz��J���tS<ƴ��k����R�t�1Q6�2��z�jĭ�fT�d[��Șj�b��"Q.��Y�:������� ���ވY�Y���F1��ҿ��b���gWwe#6SJ�cV��-d�ާ3y����%�4��[i�lX�өMD�xQ�lS�<gZ����)��E@I��*����	�>�`Mo��*wz衪�S����g>�`�������^����/|�pv�����ǆ����j��;�R���A������.��}�{����>��k��b綀��WN�>QL�LkSL����=�����}[	*s'N>V����%�1<P�r��0��l7�l��o�3�.ޓ��e&�U�H����B���>�qS&N�<=����(�����a)���n
��I)]lx%z��X�F��'Y�]]=Y�l��t���H��O���*��Zx,���3��G�v��
o������i1�q!2���EV��S�ɳo�!ܖ6 �VF�.����$kҊs�B���F���	*�S��S��J���|�5�:�8����>��컟�n�3Ir!|S��^�Χ�5�-.7%_�tV"�����|�wg����yN�>�y睵��ƛ�S#�Ǘ��*�iO{F���;�|h8P�W8o��o��z�~�^l��mӱ5&�:V���?����w?�h��OzY���0�t䆚�����\p�n8�	y����^�&��Kʅ��~)0���C~��ǆ��W�Z�3?��´��i�ǆ;�s8u�԰�/� 1�Y��-�^mƒnM2c`L�`����U1��g�v����dH�9I��$��K_2�쥟8�IV������m�҅��h�!`N����gO�4�7�J����|�/��Sgn��yW'��`
���c2�M�O9]*H/���2����.u��}D����Y\��AI
?���q#L���X]��5asۭwd��=��T���bq���RU�?�̙S��q;��p+�"�9w���$�:i���f2O��PT+xbb����n���9|�wwԧ#Uz7zV�O�M@���I��#s��2�����
ZB b#�"����b�����~��|8��L�F�=�����с�y�~�
?���E|:"�4���0�3�۲�s�*�y�`{�b�0	��g�df<KQi0���^[?Q:���_;<��G�,M��A�����
�r�b>3��L'�_L�B �:73_y{��j��ܳ`·���Uo��M��̴"��7�T������9�	s^H=��L�K�������?y���[���Yׯ!�z뭥_����5�u�u�Z5e�e�|��B��p�L5���� q�\[�0�5�'3�R_*����U��\z�'N��i�c�@���p��7�a��8Y���M�&&2�N~��O�˗	����Gؔ�z�{j���}u�C
&!I� I�id�� h3�����vt��<���ܘD���F��d�0dC`�+�8yr;�a��(}/�l��
.Fb�o�Yg����K�=�k`��w?>�|��B�z����s�f(��ԏT�ٳg�T
s�O���~�=��c�d0����Ԭ���յ0��Rl�Yf�05�y��ß��ñ>Tyr�GT���OD�&�KÝ�5[H�������^u�!%�L"Tc��v2,��m���a��c�c,�y�*377�0<����>������|K��&��L�W�w��a��2��c��58 3:����ܡ���L$��f,2Q7W�Ŭ���O��O6S�0��Ӳ˙�<�S��f����_��V��=q�^�����B����Ioq�'b��$��*L��Ku�Z�g�DT�)]1�kS=�L/�"�B�1&U�1'!쾬�DdV L�����՘�$x�Ɋ ����������X����E�5d��a
�D�+K�	����S78 �r���b�L��iې��Vd��'C^������r[�Nx��fq���A���ΕݚiV.?��psq9k #,8�	ǎ+�'�-q3)$?*��oU��.u�3p����'�����	�(��⻸,7`�&���F���1�vUN����S[f��?���/^<�>�53a�0r�~Uwڐ���|w}i��=t��0����������
!,�N<^����ʦ?�]=z$��ܼu�����~w��x]嫬�GW���S�����t�✄�{�J�3M�%	�2��0K����h��9q�������VT��M��3l�$]��f:��8�pC,� �<u���O�����	ʜ���!]cYy�Ր�"=S�����P�'X1�c�Ϥ�2HSf�}�3xNc=x�p5v3��F�iu����6���s�:��n�%>�Hp���Y��[�{�bNHH#W>:����Jo���*��2���䙛�W?+�>R�.涅���r�^�VP�� P8)֥���NLGVo?��O����Z�S�.� K7'YI)W�R&��1"�=�<�NBC�r��Cplj�lka�!T9�0�U<��}������M�THM�N8�����1��+���"�y~^�Z�"�M`�><���C�c�b۾AY�Y�M�M�I�;����&❧̩H��b-��9H�KM+c0�:�^������}	��|�����{��b4�o���LV5S���͜QC��Ou1w�̰�ṉ覎v4���{���C<���������=�2��~�a�������]����b�7Gv_<���@���j xf��G��Y�2vlf�w����^�BI�t���|����0�9�WQ�^��7{��/�[/�N�,8	]��g�6������E7�0G^���������V�X���%SFc�ѻ�DP��`^�k�>4.�����Rl��PK�OT_\��zZ	&����~G� ~���a�e�&��'��_��:j `0}�`R8kj�P=���^���翨����_��eW*+_���>�V>��\,A�(���E���ތ!�1/F孨�幩���6�s=v�ԯ��l��<kϓ4ДcH��Z�����\ a��U�<�q����O�8\s=zr��Cޯ�|d���X��u~f�>���0]�u���t*����}1E�I:�F��W��R轅|1%D����`�����.+�4�7��ߟ��%/yI�ʚ�f��^�3y������/���_�6�� 9ԃٽI�b�b����YPV�O�=O:0��l����Ņ���ȏ=�h��ʛ���{���(�U0��$�;���b��0����\$��}����V>�Y��A<�`�)1k*�L�p���5B��exzWw����m=�ͷ�:|𡇇W}ŗ-^��7V>�}񈑣�\�9�����<]s�&_,^ԁ��*e&Np)BE�DBc:8S�*ݺ�6���xf�N�j�'�"�H��$�쳚:̼�U���n!p1�w�nÌh�]#{�A�Z#�I|���_��@��w����z�ɟ�ɕO�@@�ӹ��2��ꩧ�^Μ8Y�l��d�88���f�FIKRo������E�^��G]����G�_
�F��t�r�fq���Ï{�[|²4:7fꖝ?���n����?���q%�)x�F{o$�Ñ�}�,�/Ʈk���tڢ�F�h\wá���_�=�|;��o&q�LzDuRi5���AF|{|ː*�t�1�4�F�c��b�cY�s��O����bHa.@���d��Fæ�U�W��K�U\����ڥ b4LAo�������ݧt�G�g���f��L�]�|L���e�|����<z\���`\�O~�X��&��V����Itp=�YϪ<xIH�/3Qp	w���;+ǽ�� ��]/�������T<��m���o��o��"8�f�/�@�s���7ɣ�r���{۱y/�G|���׷����;
�˼����H��pUpnց�����.%��RI�{��jW��������piĺū�@*���\'$�"q!B0;FAqUA߼��P� ��!A����xؚ/��aqC��cV�>�"6�)��\��������m��1I�$�;1KF^E5��I�ybd0��� a
���l 	�Sy��lM��D��q��b�^����|����/oD�_ǗzHיJcg�aF�wy��3���wS3��~���C��O�W�C����|�(̽g���+����NX��Q�$`#@�O�~��pU�<���:ea'�M�iѓO���p]�[�ssM�Z����R � ��š{A�{��'���Ge�w���U� 2奭HG�b�*?i<K��}^�꾥GX����퓢�NT��y'/��8|򐯺�/o�XC�W7���=�I�����m8j�>l^��Ă!O����,Nz�p ����\BY\�+��dA�^�Ա�ȇ����~�d���p�'��W/:�{0�]\�$���w�������#�F6��$��D<K����ٕl*㣒��~�n枞ܳBʙ�:x�@DBE��0�4��j��qk��@*���a'�	f�*KM�T�X\�e|�ffS>��Uq��)��y�-e�����
LZ`w/�l����IR��R�}�O�W6b�N��ʛXjvh������V6��[�:&��K>�3���w��3\��[�n�!���Jg6�@�����\z(*ޅKm���R	�0+�EP�^�p��}���7�T�h
�u�my�$wT2��+�oG�c����l�ds����Ԗ-��L�GՉ ��}7����B�]v㬅�?L%ﺙ;��A�M*kUղ�PHѢ1t�g>�9�'}�'U7D�k�dIX��b&?�c@f�)��o��o�Al��=��YX
8"�f���ַ2�M5k��;ߥ���㝠���it1V�&�|G������`$!)���Oy�]]2X�Ay���3��g�E˳M^�W���Yj �I孭���`J\��:q��W[l*�:;�L��H�����{S�ʿU��-l�4�u'ܔ)�{��N�i������|Wwxڌ��_TO���V>���]Y�X�Ѷ	���?���6�XP���~���mA-&aM�k��(��1{]�T�p�D��>*ܙC~;;�X-�t��Dب�،-z@8:,�ihn���1�]̔9	a1�[H���������Ǉ����wv�W��6-i�ک)�V�Dz!�ɓ���
�w/�Ęm9����F����KM�PW�~0%��zw.�򭺏��덾w�]́CL���1R����@wT���27��_�,��C��y���9e��Jởr��d~��ձ�%�y���3ñ��m�V0ƹ�Y�p�    IDATtq�E�[Io2��g"������DE����Z;u~�;D��C�tԃ��B_  A�tT�k�g|�gTe�O� l������&����@=���]�3�X����x��|�^��1-��@1���>M���ǤHغ`�p��>'�tZu��ީS�)���
�3��OY��{
i���k�]����MYʁg��h�SO���x�[���o��֞�C���ys�M��mo�����&��� .���{�a[Yd`������pZ��Qm=�7���X��wzo����%w��c��`�T̢p�X�Ŭ|���l;�=��k_��2O5�Dwm*�Jw�v�L��A�!D@Jy�ePF��C�b֡1'k ����-�p����7���n$g:�N� n����� b ��4&=�qkWV�	�p��y���ş�3�̅���Fm�6&�Z���@�Q�J�gp#��˦�� ~y�C��5ƄRW#�D]0��0K�C��&T����y��G8�=F���i"�L��S��z�%DF�tu�'8��5�&�¨�6N[�	q-��ؕ &���튛�U��&�o���%yL��[��$�Ǐ��-_�0U�	!��Co���AtSMvK�
	�G�����OG�4ߕԇiH̋ M�kcn��ʦ�RH�4�"*�aj�9?U'��4�λ�1R���a4V�w������\fW`x�N��d���*����3��{��Ge	��=�z�y�'��i��Q���]���=�Й<��"5�Ӱ|�HZ.z0x���3���k�N�h�<�盲HO�~����W�Hs���6�,��7X�0}`�Ѻ�wfӝ�����~��p#dv�\�6������^�Ե�eTN�rl�fT�������'Δ]���bOv�Bx1�R�H����2<�݉�*�Ņ�u�͍9�s9��>��>$5G��3a�������;O�ܔ��V�Ӹb	����|n1z�v$H�Do_�
3MD�υq�3���Ҫ��w�b�*ͬ9�}���po�b�����-/ݜ�"&e�հS�]l�N��l=B�Pl�f�Y0̠S���~�������`�Č؊:d��a2�;����0��fEL~���7���a��N�������`�.�g�ٔ�8��l��R����q�8��̩�l� ��x4n���HW{��/d�k�F������Mo��o$co��>4���?��GR����lK���L�"�H��R�)�H�npk���嬄��B�����[��i��Pҵէ�9>��8��"�쇇&^>��G�&��,�!i!���V�֟��Mri�Z&����Z�����F�)�߿�67S.��8̍�+�Q!��NV�H/_�%(�3���9�I���H(� +EF	׶\$O�ϑ,8eq�$��J�Eˋ�3�"7�v�ӳ�<;��t|];�-�8{��HJ6��V���y*`U��R��A*���3���
|�j����r���,�=w}cex�3��_V�\<W�� y+S��b�V�=:}t�>&��=�sa�H��������)K�Ƽ��v�ܩ�jȔ��JJ��e*����u.��_V@�id��h&W=��Ne@I��c���9����@ʣ�{��ѹ�{��H������f�z(��?H�?\/W�R9KU��S� �!�F���=�����ѧ���Q7���m���b���_�j�H%�Ę&u� f)��u��?�Aˁ}\U�{�Y�ɔ�N��EB��J��H-Ʀ�|�me�Y[��1GE���b�\٬|''V�^�g0�6Mn�Xوq!V��Y�Y*@V������]ԣZd�!n�����:�;��f���CK�5���~6W�~���b����9�6��x.���d��?�W�7�t} T7�=Aؼ���Yw&�s`x��4��e�赳�fz���Y����l|y���ИW��pg�w>4�K���2� wzo���=�3LM-��9�{���|�~=�v2��O��������CZ����a�ލ ��
���5���g4NZ�	<��q���.w������/�/rH��u��Ȉ�F�=Db|2�x�U�w��rq1��L��ed��^��Ft&D��K.�dƴI��ߎ��3�E�u���I��ﺷ�˂i
��)y$ݷ�51���
�z�ɤ�SҒi�nX����ұ��xs<�߅0��ӏş�Ψ"���I`��
���G������Q� v/0��RlõΞS�-&̪&��=qӊf'k��ѧ�����Q�Dz�Y"øi:��	�R�4�������۲��7.~YH��x������O�F!��=��͹���^?sOd,c"�*љ
��r6���~����mk��l}{`1�	�=xv2Q>:�=�����k2-�:���0� #(_Pfop���HI��@���4���a��mne����t��?�>s����ax�;ޞn�^})=J,9�g7���3y�wbVz�K��P����I�+G�ə0VtPD�@��&]0\5�FOc�ы��@=㖭����s�3֘�}���X�Ƕ����$��]	zШ�a\� �@Ofܠ+tf�X����gQ�,�)t��{"���3�bf��H���8r|������S��o"�e	�����L&C��/�˧��؊��L�;s�ԥv�M���wT_��9�+@()i� P�u�C�F] ��j����./>0�Kr4>�����~c|��L�o�?��h���6<r��4��OR�Z�Vq倥36��,
�6XL����</^��i�s��������E%��r�+�gx��o�r�����F;YW9��#�2��������i&:����$sr˗����0�D5x�4+�2pԣY�y˭7�w�T����ca�>g�!��,ڥ����o�:�K��q�ʇ�Vf�4F���Zޙ�G?��;�Q�0	�{�k�Yaz�jzF��O�e8�	����vr�S�>;���s��إ3�1�Mdq���[����h	�R%m���ۓί'�O�/�G�u>�#��ѹ�����~t8�K��f�T'���R�ŀK٤e%��\*�E��]�����GO�S�}0*E���d͆9����{�D������".y"b�ЧtK�tx�@��I
#�6�� ��/=��lu��t���><��E�=~��񙅽s+K7<����qx�����v��n�	j{`k�o���������6]c���$4;�r16ɮ�!�3V/�������v����h3�5�Lfm�Dc��>�y�3��{�}-�w�+�̰C�97U�0N��a[ωR��=��F��e�͑M�~�'~������Xh���SqZ�f�'��>t��`9��U֨g�	�24,o���ն�����R5yAR}�ę6��-}#�/�~��X��0\�Zd�>�c+N�Y�ވ�~$��	Y�#$�hV�<ЛuM�#=�h[Ic�IȽ+�Ҟ��g�$u�R������p����|��F�R7Ds���Ƞ��T����y&a���t�`y����3x�i�$Ji
m�Ù����Φ+����ٽ3{�9wr���S�-��4��7�r��I򪃺��#r1Ts��}ߌz��7����1��O8�RQi�nW����2���'>e�=)n+����'����ު{I���Pp/�ш0�F�7{���ѯ2��Vgz3�S!�3مц�`)�V���r���s��Cs1�M�ʼ�������G���<s�Ԥ��3��6����#ێ���d��YK�Ӷԁ>p7c�ë�N�����c�{����f�">�����̗��\->�U��!�$�.2��
Bd���䱱�NY����}�Y�[����k'O��̆/��A{h�-R3�ɟoFR6��K��*�_��e��7�DX�Wc��㫑�����Z]����H�Ŵq!��}ss�1�/�LxaJ̠q�I��^���������~�NoC�JRS�����=9*�9�l,�ؿϞ9�squ*�'�28���icnj���ō�?p�o}k&B�H8���p15�Lo�5&7���z"�z�7���F�+��YF��4�e��2p�{ە��?�����K۟��>�'N<~8{�L�p�fj���n�p���Bή�>���GP4̠9��Wd�2���O��g`xE�k��f�9gH�j�1� yl��mE�9���G�sf4"_�����k���Z��	 a��)h�����	�����%�r�Y��)*jCt�c��0�!�gG?/�-,��ܾ�ӳ7�tˑ�CSQO�]f<HBL���<I�����2#���ZE�q6���w��$�%P��e	J_��'Oon�.-�lLL�Lf����ٹ��{������x��K*v\����t�Hs�2i�z�Dj�SzyI�H'�6`�7ͼ)�9wv}n{ϙ�3�1�������'w�N�n�D�����֞L�M��H
k�;�'���C���춘C�G*�l7���>&���+��]��̧�΅�&�{�o,��ؙ�Iٿmfyssgn+�O�XTM��0&-���d�2:���@�����Yi�.i6ih`�j�>뛗67���OrOl���g��������z�0MB��*u�,��X0�k�tS*�XEUx2�h]8��mtm�<4����,q#߶S�����w��C�fl�v�"1�.E�f�)/���P��U.�8A
e��6��t��0���T~f�2�����p�m���^��mN�m�Y?������d�:рL�'�1S�HP'x���`���tpfѭt�'�4L���0?+�U"xY�Z߼0�x`}'{O�]�ܘ�[����{�칋w�F߿�HA��z���5��&s0�F�lF
ܙ����D��M=���5�g;��&h+Ri���Vv��$��wi�dTǙ����'�/\���[/��l��,]�w��W�^+p���|VU�����1��3���qqq��㦓S�B���$�'����8����!�y�����`y|C�J���&D�����6��:S�p���M�ܺ���?k�#7]���_��޳y��O;��Ox~I|]�AZ�!䍉����m��	�����nNC@t0�8q���F3"�b��{��ژ|���΃�k;��V'Xߞ|8��^HCٱ�K��h�=�<�ԙ�;��x,��ݲ�l�A=~_��QA6�m��>�|~����2�����(��֧c�����/�용��sv�
>���-Ѕ<���ԡ�Ϣ>.?���]:��V�������KS{�]�
+��{��ت�9(K|�k�)�\Fw�v�#�\�b`h�Z9�H��W�6�� ���������}��-��0�}�5�K���!� ���������`Ez��fPi^����)�߰6�pxmz����ҁ�#�=���LMo����̜��B"�� {|L�!)��HF��b�R>�$���\�'\^�=��6������k'�6���{b~~��lTp`F�s�i7���z����I���3��&�U����yHc��u�ңŤ~a��օ����m=�j<x!������޽ϲM[��V�0S�f�+�1X���%e4����ϺJ�Jo��?*�Y:LP�� ���,e��g�7^��l"�ށr#s��[ۓ���Μ���3�͚�� Rwu�wM��'p"�$*A���i&-�E�d���I=��'��\��/�NI `p��жPݲ����&4$v�7�}]%�?��U$��p�\Xv>�=��V���,�GzڰᔣA�À���ș�C4pv&��Q������յp���nz�͜��_�ޞ٘��<�g��b�&Y�fg�lӋ�����5fV6GT0�jp5PJ#�p�+���tM����9Vzeckw{*:mN$Y���z$��F�S�/�L�xF\f4S�2<c� ��Z(�,G|��l��	&[����z����<�F m��~��]nw6�?���/��5җ�VT#�*���p��P�{�\�C;0g�"O�k� �5�c��+�.�6��[�%�I;Ƃ�w�=�xf����uUwC�4q\uO2sy�wn��n����͘��Pj6JyVi�>��\V��:5�!F!:� ��w��t�9�C�Mg �j�L�ą�.]��{�衻�3K�w&��9usb{����|���}WO�>���ѣk$����:B���O�~�zf�^����2�8�0O]#ť�PrIqM�]�ڝ�>�y��I[�]�!�s;��/d�l�`^j�C9�u�QM��P���x�iO�k��o��{�ynImh��ɴ�)���{k	O����}γm|��ęǟ����s��#/\�p��˧�w��cύJ��^�o�:���4��^������z `�<��5��iqa�̥���q'��AO��Z�鹷����_����s�V^F�|���F��ٔU���~�g�$�V����񇫲��K�]��m����;9�";�nf�y��w�Ο={0�*�:}j>��5�������)�H��#S�����a��k����،����F��_�ar��-7�\�V��.̬onN���w{hyl����e�S�졝��ǚ2��w�k.<��&m����w�1r]�}�;w��{���7)R�$S�]S�,)N�q�T�0M�p[@MӨ�?-�4(� h�(��H[5i���Ӱv�(�r�Rd�R���II+r�%�=�;s���s�^�bH�"��V�^i8����������A��kQf�@|6�駟NLN�H���|����f�TX|Y��<s]ŚpŶ�:�-j���R�r��6�7��di���ā��X#z�R�R�<Qh&����hK	f��{����}��g�]�w�L�<��(+�1Y����Ɓl~�c�-{����6�0a�z�x���M�5k���$"�S��㮻�2 ���W�b�
p����#��J8lZ�	�?R��[��`M!{43x�?w��333�v*[�����Lk
JP�e�f$3.�� �۶�+�T}�≉Y&+*A�e�-*�yQ1?=s�Tz���>2L1u�������u�ًsBL�m�`mRb�ǶL�vY���2�9dâ�s�,�����%m�R��._�|��E�2�׼��{�'ƚ��.z��۽�C�VUe��m��s���FǶ����d��������Ǹ�ey�Ȫ�Jg�)��#O��_K��ֱl��N��.�:h�����.-�	{0~ Š�r�};�O�.�-"�^��蔇�ؘ�V{ep��6Zu�-	��	������tqr����?��W��+ SX�_�N�W�.'��8pŲ�d�.����ժ����x��iYX$Fh�iwmɲ�Rc _��2
��z��:l�h]Qq��H-5ț�\v�=?��x饗_���6�7�F���o��9�%���w��O��jd/�l�8}��#�ꝼ��٩;v�=}���f�C����"W�쌡ZP3dbX�7*Vν8���[��8�de�:yR ��w���I�ڔN�.��fd�IcWd~� ��S���g����QˊmB@�����|�TP�P��*�R�R��vT��qT|'_�9�e��G����<s��lO�K�U�v���Vl��^����?��ta�B�M��{`!��}(7A�
C���(�j�mݚ�0}:�Ƨ�)�Zd�K�ۍv�z=){��gX:mUJ���7ҟ�X��X/���Û��2���ވ�;�i�-�	����+`	D�g��R��'�k�&��ʘ��X_�M2��@Q�e���*�,��X�d��̅}A��r���7ҹ�����z�����}�*�����?���c�^�3&��xO��.,�*��v�#�`�>\D�  �l�Vm(�� ��P�h[����/��WYJ$��l��BJY�8�@ 2?��(�  @f����I���Hjm�<��c^��.y���pə�T/m��=��� "��X[Pt�X�i�)Bn�FQ
�����AQ�oY#�g>��9�W�YW����K�)9dp�P,�N6����;�n��Gg���Q��    IDAT�JF��ܸ"d��������|簢7˦�{�>�U�wH���Fkc��9�C��_d�����p{�7����E��r9������l�zǏ�,�?�䟵Bnco����{�wpq�U� �H��2?iU������w ,@ @E��+5a������}�8wN�r�8 @3��4����b��k��`L�� �g��Ŧ�)<�Hy��/�ӣ���G�w����.^��k�Zbt �k5Ŗ6��6D\�ܓ{�"K���8
�N�I�p@0� ��.s�C��4�N�h��rgK)i�L��Rٿ��=��xr�9�֥�Sw%J��c۶ٱ�b�8�I'�6Wl;۶;�����~é˺����c��f<����p�+Nx�
m�ѽ����(�6�Qz=��^\(DE�$�(�EB�;hL d}~��o:�x�_�X��������`��`3�O����6�H���f�k�3s�;�p)��i�{��#+��t��9Nw���YQ9H��v�J[� H��}3#J�󹴘�0to�$H^غuQ���6Z8d�����`�Lt��{*T��te�˱��	�}zuzЛh�N�y�<!��m&[���A���J�%�&��
�	a]��.M�#;LD�~^�]�=�y�jZ�lo��쩩����cJ���M�_%��x���ux��P������a��"�p��T=�(wϤ�n~=i�u�`u�`�NJ��/
��؁[�x��$�}�aa;yU��Rb��5����9Am�{]��Sf{]tI�b�� �{����ų�����$^_yC���f��UC���2�������:j��M�@Mp���̄�rɍ$9�IQ��xrp���tUP��G�PTU�VF�'��r��d(�!�p`�q�2bH�9CV�!x�.���Z$�AA1����L*�<(|Zb�>�)�X���:�F���җW�*�.��WBW� n�ƹ�7Kg�׆C��A�%X� �p7ZLL�Ʋ.�97jz6mjdit҆��u�����n~`~�P�������Р�g=O�p� }�3�ub��#��m�1�,x�M)��M��
�b���1y�
ղI�G7�L��.\�f3���SNJw�s#%��2o.��P���^��1P	�l�֩���Y�(�^w7�#�֕F$�_ή$N��{�R�.�T�J̠I;�x��y�եlſ9�5�j�������;����0�%B�zh��f����|�K�7M��jH6Y�Y"�XG�#ѹ?�ތy��D�
�e�k�����S�A4�J�)BeQf��z�!����������4�1X�کzB�g��\����-d��a	H�G�@�8u;������OHi<G���B�?V����6��D/GQ%|�	�*]N��P,j!�D��f��/r�1�鹚�;$�aa�nا��� ���t�C�����<@��a� ���ǔ�����D�xvv��K�b�����>��
�\-��4\��5������ {C�!�D�Q=B�W	�T:2QD��o����o�[O=�({+ǲ��k�~.�x�ƣ~����f��V2�`@��7�l��%������s(��z���n�.0�ٝ<�+��״�=`\��W�57?����%�e�l4S���~0"��ZX̜77F >��BOb.75���]��{���T��~UhVFq�d�R t֑�)�*3��c�U��0��uQdE���1��ڵ/�C� �IU#�gg*A#��K�� �-?V�L�&�5�"�2P�D��X˟6u��.s^�"5\[شS~���_���Rb���,H�fT,�`���!�x�O3Iw����Gr6�3$8|��D������`�!�N̏�(�������n6{2���J���!5S!NOh�Ta-��o����u�������
��[X��?۸�~啖 �k�[2i<P�̂V��<G��K��É5���FHǲ>&Q���u0�G�BE���X��Ua�f5��#|������}��Pa� �n�}�/�u|�2��[\t��O9&O&�+Lhd���rH��\���'�AX���n�k�5ĆB���g2M�[~� �a�qy��.c�����A g���������̉q��^?	�.oYBe#�O^0��_8�m7ܗ��ۦ���K53-^2�`��$1�M���M�w��\ψ����qect�䝤�i��}۳�@��r��ي��c/��C�/���o���n��5�\hТm8C��A&2i���tEi"���ʠ%���>��b��~6H�`@����.y�ة�d�n�<B{�攊9��Hb�@iS��C)�l���R���Ur����a�{B�ru�����K�H�0�*띃;<���۩���K�o�6َa�8�I�[����/����y����B���y;����QOM�t8�i��/I?k6�K�BXb�$Q�զ����tb�
]
�)���Z3>8�6�o�aV/�Ŋf���2kB�Æ�c��k|��մ,ސwR��$
���<�l���M^���cS��)�t�㎛g.�!D��o4�-m�%�!�d˃v0v�X�v},��1H��1!1uN{���>G�tz|Zp��<4�ۤ�t˞h�(�;�J��P�&>�F���1��m4�$l��2M�%�)��*J���\�&^˱��*Tk
"&Eޙ%L���u`z�;j�����	��SFQ��ˌ=XK�b��������2XM�a���$5!�jd!�Y��0	�jޓ���>�������J��W��;���7TD7����!���������P.��f���T�(ϷE}��t^�>C�����zG�pȭ���z��/�_4\s�R�hqD�,���A�ɞ�(���-뙨�����0�0&e�2���a�P��Ź*�dQJfy����_
z{�)�z) ���=V�+���U�Q(��Tsّ=\����ƂsLP� ��%�Bq't�Y���|�q���6��|���o2�.l ��ńQ��V���`��޳"3:�p�m�W�m��%_h�x�����xB�H}�ėT)`��r�2��wD��a�5z-��W����-��mG��YM5*���Gbd�zA�����JU]���C�c7����;ClXV��͎��6_�+�n��[�A��l涡$mh��6e�v�|*,��::��\��`+�|[��R����:d��Tn8�"�?B�#SddZA�^A*�( Xp��rQEv`���5�2 dBt��"�w�.:b�8(#�m/8�E�
M�H#G����I���*�b�� �(�^nͭ/-�(����yR	 ?�yҝ>��Q?�w����B�I187:�e�>���mE3 S Z��k K�2`��k��p�akBI��1�k����EVmO�\#gO�/��83��͇�a���m8I�y�̔�.���Ի�'�d����8��5̣�0S�ծ�������Ξ�Dz��v����ʽ�	Kus+�Aq�'',�Jbp\!e���i�W^J��(��ӦI�ע�F��4��9+��F
aO�jQ7��W!��:�yf�$i�S�πQ��2�Y��hk���U�QY��A�����6[y-����0Y�^ngK��<�G�+
+%N�a/�w�)O����fՂ�L��*����G��>%)>�V�ƆjFm�o@���˱��'�j�є�t8������A�z���]�-q�L*Ng$���@J���y�3-���l��pD�e������Q��CiӲ�C�9�W`'��l���y�-r�����2hEa ��|��6v|�S��tU�-���uܢ���v�U9��H�hP�7�4B��1t�(̈`��.�I>���ݶ5�x�2�w�ni�<��`T�vғE�TSi'�;�2��1r���uS�S\�.r4�R�~��+GA2����@����ܽ�2`�����v�R��'T6�β�[�:⻪�x��BN*@g��Q�|:���Cd$�w#l�zC��n�������Ae��D��(����$b����	�&5��*ϋ[-&CK�W^%Ï4�-�a�0�^��`���d (�MON�;�n��6���ޯk�Φ�U^C@��q��2s�2��7s�;'�#֒�܂���|��|đ����ոu���u�Xb��i�+}]e�=B�Ș7�H�)|���*���S��=�oz��~rdr��kkUo���TJ����T_�1�d��M5�Ũ��ͷ���$�`ձNg��xz��!p��U��,�Q�v^Fr=Re�%-��G�]Z��/kguX����=��'�����e��U��9y��u�)���	pQ�Z��L�0��tt=lo$�[�ʳ�;����`=l=���f�jX�aOHՇϓ"Bb�z���w�[R~3}'�NvL^QjMf��lD�Ɗ
��Ϣ��r�4�i��}�d�`�r��~a��U��)��V9�i�qy�5�R=R�+q�ɻ�ʹߠaW�)̙Ħ�{�W�H���	���\q�3�K��~n�E��-2����:[�H_1Dוt����������"�ܥC�ʪ�[���.H;��x͵���$�����;d3��u'�rhA�;+mwtO9Kj�F#_�b'�/�dN��X�m.JK�B�Ѧ�[�]]qM����]�1��̷���8*����oᯀ��7���lT%>	��1m���V�%��y�&������"m<>ː�Ȕ�!~�ȷ=�����+��
w�D�����KZ����6l@�F&%�4��N�J���T��b?��ߏ���Z�J;�wۢg�+�D�7�U�%BN�7hg"�и�իfXݲ�����x�EC+�}����sK��(S��N?���߽�p
+��%�x߰��ˇ>I���Ŭ�΋GE���{y�.�'�'����v��g;����R~-�9�Ju���@ֈG�&��] ��q�I�[���Pǡՙ%t��j�0�'n�W�cK}U�.�06�PwT�ڽky�5�O�+^��TMϖ�Ï^w�Nl@�ɾ^�j?����<Q����*�8Sã���~��d��c��;��M�������G5����r�p�ͬ}��~�~�Ԟ�z����3e�spF�Jmz����')בd�Zʒ�@��Ƌ�s�d:!�/��5�}��g����nvH������;�	�n
9����e��bڴ����#M6(a��K�F��{BJ"������T����bn0���a�[�M�仝���f\eemI��K��p� ��Q �³P-BKfL�B	Zÿ ٲ���8;�]2�m;W��n\K�RQY_�R"�p�Jy�w5��(���F�+WO|�5\r��1���l�E�Y2���^܇�`�F��ʠ2�:a�/��jR��m�T-�cV�(�@�Ռ�s�������f�C�_�"-�a���.������J�'�Q�MԴf�<hPS �W�P�ǧ���O��v�^}���J;.-�>��G�y���Y�H�{��#o��3�D��ɫة̫F�6)��$����*�vuT��j����5$f�5C33�&;󚙝�)R~HA!�'cf0I˨�J�ȔT�����v�o���x �@�YHa��f����.�O������k���<���L�,N��l��lI���j�>l��*���.���	�� ����0��Ի����C�6:��ki>�"��ע�[cCM0Aň�6�`�,��Mm��D�dx�K$M��&d�*E�w]K�K޹"yL��5n[ʌ��A6����+�� P���-�q�6h���4�I��ج5�'�=�&@o�U��y��DLB������;��:o7m�����o~�F�C�,�,�B
>ྌ����,�%al�e�����r��څ��?#考̯�=Ws����d����%�BO�_�OM��ë���K��6�����5兓�$�Y��_�c���;S2Ȱ4�7�s�/ȣ���IS���dx/d���v�H��R�H�F^���0V��ȏ�w`M����cF�`Y�C��\n>y����>j�,¼��8X4�QE�Cĥ8֛H;WZ	?I!@~x�8��F\�\M]u��`]T�o;P:�0��yE�d���|rĘ�� ��_��]40]\���.�ktO1,��, ����k/P1@�m��:�K�`
Ҁ��B��
M��b3|�v��,���΋���4�D!��F!|����6�pza\�%E���l�i�$U8D�Kϥ*���<d��Ҩ���nD-aRwE�.7aƏp�����{Z~8P_�ľ��N���B�b��品�B���a���L���ז�(�s-n�aK`��B���8j<E��Z���בJ	������	�%��﭂U�u�<�|?�bz�#��v�?>r����MA���[~;�K�
�m�p��3a�k�̬*6���l�oJW�n���=:;Ҵ�p�Hb�5�kw3?�U���ዳ�$��7�M�j'�q���vȚ��Ӧ�#Zz3>�L���$
��
�[��&7��E$��鐺ο�1����̠��b�����]\��'Us��/�ش3�DM���4�_m�M1��*� Qw~g����n{��ɪ�y���Ǚ��u�L�҄ȣ�G��Sn,5ÚX�s�_�r�dbmӗ:�x�6������'~+����Г���LU�.]�{Ԉ����h����j@����'�.y��x~�	_����MAsñ�6�<�o.�??+���Z� l����l/��R 
_�1.��x��ݤ��bVM,��Ҧ�} {�yi����+w-J:��'ko�|��#i,�j�8���qfhn��h�ٓ�Ԭ�{�a@B� �F�e
6Y Y��̷W�^��~�R3��St�M�Ɇ	z}�jw�aG[	_0+O����@0I��ק��Co-��X$ĵó�G�������?���d�"5�R�3�1�����ӑ�@��Y(��j�'4��	����@3(^bܕt��'qC��K�c�EI�Fn�����q;t��J(�t��N�ǭAO�$��JRO��'<^�!mXL����q�e���(�Q*�]�1��tC)�{QY[��y�M�/9�|*�t�QF����'��!fl�VK�zS�'�fE^�)(-�S*���q{H��`i��=�e&��֙I��l2q�zT5!���.l���@�	��޻n��&�O��1$�[z��=h|`̒��n�%�����7�,o�:V�ыB�
լA�`�aW=AZ�$���X���B���=`���F㚜Z	��T�i4�:vX'���!�R
����<;"�_�+n}�a��AE ��5��t?D��5��4'\��K3ɋ�M�a���y4O d���J��j��$nǌD�g�E��)��"�
.i��1��ޟ�Y(\����I�R����v�a�˞���x��TΥ&��`��
7w�g��-���y]h��1;�p���F���\K~���&(U&�<ᴤ����\���C�Hװ���4�	��d�Ȅ'����U���*�]�`j�
l������5��IhX��G/܄r�7>������Aoul�v�3��<�% � �:j�:����F5Kq)Bsc
zbڤ_���5ɗ� Ե0Y>��)�T�<P��gX��;��0K`2�]�����!��:��7A����`�,Y�A=���W"nC'53��,{�Ȓ�lD�F� Ib<OHA��tk����pܪ�wL����:�k����a4�K�`I�i]���v����E�'�Ze�@]�V9=�����dzB�H���g.�B��S��QU�+��Y9�9������Y�NR��t)=�C��
1�$�@6���/f�&hݼ� �̻C_�`mȏ�|�}�+��j
�d��&&~��V�]���]�/s6�S�f�<K�$s��Uڲ��sJ���0���C�P��̞J��|��2)�y u}s܀S����c�X܅G_}���O���y�<Q!��,-��?bgo��Y;������ []�gw����0�tĴ���Z�d�d�O�O��uQC/8�՛MN~���S����QW�X"�D�'��	ٵ.9���%��Xs�����/�Nw]�L��n����my���v�;dCF��C�M�1X�	%8�}�*&L��7�g �4�4�Yc�b�J�8�����^f&�vz��>�4�(��İ�|�	�@���Ƭ[�2�.�9��/�<��*n.���f��%Tg{8��I��.��D�c!�A�PRM��j�<�T�_�A��fG��U�*T�;l -�/-��*k��K9P�����^��j`*b��iv��IbAr*��y>aƘ�
5+� �sW��6W��	�7���^?�I/���}"ژ��.V|<:!+7.���r���^��Rk��j�02F?0���&��*�1�5�\&]]�+�|�' �\}^"\���C����
��oҚp"ꀆ`�K�(�7%O�a��l�����հ>64A��&��l��ee9q�G^���W��;�us?l�ɥ��1;-,S<���)���A���z���s:�f�1��?G� zd�O��6Ć4��zֽh���a0URVn6�И2�9��_��{)R,f�e=l�/���#����ل�����ʊvȂm��Ts�=Oz��B
���Ȑl�P�,���*��,DN*ZU5Q��>�:bXj�e��:O6O���
�|�J�6 L�,أ���GkϾZ�5�^\س��j�xi4x�aA>�T�zE��)6�&������%u��oy߽�ч������wF�K~�:���}
��[��D8��7��v/������U���L�t1�3�t�KT*�.\[C5�7�g��f�:�f�-@b�k�E`A�*�sd��o��%]J"���z(���Y��+0�w?��L}�7N�����x��GI�t��^�����Xmb���	qw�� 8-�9��1��j�����e�m��xUM&?2��1�⠋Xo���LPZ���C#o4Su�Ip�?u�~mg4�qb,..�9ΗKսi�XU��7⯢xU�ē�l`�3T계�����Z��~���i'�|P�T�+j׮�c	F��u��f�4�h0�X�eb���5����3�����4_��ӵ%�\bg\�� w=g�$�������TVR���8P"��䞂,�����c�83��qU��S���PC6�2<^8�{�6�Z-��y쿦ȋ�P���1+V/P�:�}�s�������,$��TA����Ocg��s\�=��� 6H�2�E{�)S$Em�D�k2�MeY=6�Ϩ��E=r������������	���
��	AG���HF>Ӵz�u^X[ȟ:k�.:aybl�voΖ�eB�E�_�z1�(�߾iB�O�@��QCq��V�L`���rD-E�b�r[�7�t���;�ۈ�^����?��K�n&:M��� HB�-�cқ;6^�6��J�̵x�����#�,�?��?gHy��'7�c|�>X�t��6�6Vr�.��9ӊ�Fvv�ˑ��L��6&����?��s�RJ7�H��J��b@�Lqf({��֨}Z�����{�@`Q�u�)��y(#A�n�����6��1�ы}cd	�!�	\]?�ǹ���'� -'��G�j�}DpM��P3ETw���x������^}�%$
J��7q�{6jQ/�b/'O��G��3֖X�꽟�����=A�j�b�! ~+�>t�
��=��l�@�`����Z��[�
3����=��4%��B>�C�C�#��Ҋc�S����э����l�*
�%��iUHu�3Z�#�7b�G�f��~��~1iA>���f"{9����V�톼o��5����>:�y)),LI����CG�֎���8�f1OO���m�&�7��G����	r���c�9�B�A�CО��w&|i񢒹ʹ��������ñ��i�闱P�d���P2h#���|�V,)��[3�����@a�2�)�������h���Â�<��zD(��D���̐H�F�X���Ԝy�T֠ՇprЎ�.��@:D��L���'g��mv����qanv��}�����
�F�^�fRi�d�\lxi1��P��+�| +�u�j��s��o��kQ��V�fR��Tjxim����f�q�&^�f� �B�JA�
�&�@��پ��ր�J��#"� (��"� �;�<��X` �؉0p�?d*@�&�LP��c�G�F1ϒ��N�i� ~���^J���n��:%�U��%o%��h�;x˔]:,g{�H �P!(�^��H
�?x���y�#%[�`�/��#�?aWuI�UY��w�͐�+BUg��TJ$,��I�ߌ�Ҋ>l�T5�C�V!\��<�z!�iw9U��/"�?�	��#��$��aK��1��4 }
�$g�۱g&�g2��B���V�"��)��j���W`X��`� ��c�$�t����I2��	�W���=�h+�41 ͹�S��B�v��A�!GeM?�s�Z�k�����Y�8�T�X=VB��9�d@�$�ԾLFυ\ycei*
^��Llbߴ�\�B/�a�5f�W�0ر�1dwi������/'�9����9��cn��%zR;M�΅���1o��i���K�XI�+25����6�Ae3V�g麕I��F;��Ѳ��J_����0�j�����5��ܺ�d;��j�`@k2	��`�֚)z����k�4�C̓T)�a30ǔT����~A�;ӵ���uϋ���Ș-|���:'{��]c7����*b����`?M*��c����9�j�w���]�B���=S�����VϱA�.4���?2�	�������2�GU��/�Y�D_g����K^7N�OO��'GQ��a��`c#��b������Z�g�l躚G�ٚeT�O?$H��f��<��GY���=����74�ۤ"��
��@��y�3Sה��q}5�[l5�K�6!j��=�����o�t��*���f;ZV9C��/���S
,�+ #�Lqc��F Y/أ�A�c̀�Z�У�n�ov�*W�El(�01�8��6� �;���l�
�ҋ*�uq��6�8Q�1a�ID��/���{c�$T7�'���0|���{@��D�0�䰉{��,�1pp�I*R�H�f�ş#�x9Y�nujab�)����6��ā{ c��_}	SR�b��Ճ ��}'�x%�H����y"���h��~��-�ZS�&�p!� !V��u�j��:�bK�*���y�7"U
5�D��}�F!��u��Z�*_mN�Jq�ke�\����|�Ċx��W����X���#	&��L�$w֩~<N��\���GL_�sZ���ǧ�s�*R�\��Ъ�e�*��:��"���Ֆt��0�;N�m!3I�j?@?v�P�H:~DK���"A���K���o�Am\���%u�j��\ދ��3�}��dq�W�U�a���X���rz~��c̠Z%�փ��i��pg�E�_0%�\p���X;ђ�.	ѱ!6�̄oɁ���~�F;0��{�D�"<�y;N�a�hF��#��}A���Ұ���r��`�ڞR���F���JǬ_�c?��'r���k�oh��`�K��델�}*�E�=��ᶨ1���|�*�iTn���$���x��#�m�������aǎ|��FH��$+�sQ3e�dХ�\���IѲ1"�?>��u)����Ĵ�6)/X 3�:���$΀򯻣����� ���8̫���N(�P��V��v����r�%�K[�m)K��b��������R �����_��������:.BmɎ��θ���i�-�y@��W�s!�7��ƀ��A5ȸݎ̙�ń�hb�4��9��4J�/,�y����-�y��z���kh��$
.��iZ�)�h�pX�5vNpV��G���x0[��7�tVj��D����/I�3�. �7H(}ͼ	,j����hx�q��OK}| #�\�l}��^�y�&G��?,�W�Sn��TU�g��	%B`���Z`��c���]|�1+C��3�8r�>iW�)=���a�?U��׉YT�r,�q1��č�k$�4�t�����ӣ���
o-�W+Q�ԉ����*C��z��&�7�qq�c���T`e�4,��zX�8������	<��\H}�7���d������0}U�&dE�����-FG	F�˩�����+�F��ؖ5:����	�����l^��NT  ��T�,cHzs��7Ե�40G�d_~�@��^�_�<��3S� �c�l D����ȹ����5om�G8x���4�� 6'��֒E��!�Ú�����Ϥ����r��'H�T�z�`5�D�?�#�S��%�U!�&%ww8�<����O������ѐDN�:��H3cd���|�&;�����C��v�Q	V��Dtl�qTd��bw�e]I���E�^�)�!Τ���.�b	��2�RҜm�r�~V���y�u��/�Ou�l,�;&|8���Ο5Rk��1tkΛ�p�*6@ƫ��y\L*��*i�%�;��������Mk��
͚dnï9im�(D4b���n[�9?W7.P��7��6��Nu% 0�G��WT'|
��p�#MW��*��X�4�BS񈉕�v:tF,���Tx#i���>�H_O��K��(�~U��g����##�a��l?�� e�g��u�y����)4�H�^��h������3NU; \��
��l��:y�D�`�����unlc���4��F�"�:Gխ��^[,��;L���(V�'1��W{_O��$���m��i�e��Z�m����Wߺ���j�L]�u+�Ꙩ��a��sZ&<��G8�6���E��?�>�;m���X�P��9�Jq��W����bH�y��HW��~�u���B^�M$I��L9LLUh�jQ������%�Z��@�/��&�[����=Su9(�A��D��q���v˩� R*��2�0`}"��V��n[w�b�i���躞�%&������<�����Ƒ��%:�OE�S�y_��|?G��{�(�ԦO¿�g�1�y��b�TIA sú�i�t\s�J�Ū¯�j�����?}C}��ǚ�}t�gÂO�un�4.M�% X�_����?�����u�2fD���LSg�8��\��.2���y�T����s�R����a����̌��/F�;3�7�Ѹ+{���#]�۶y�U!g�;�f��.�ѲK�@��[�0��H���^^>�%Ha�^��.�Y��r:�i�|b��t�ۮ�M��me��M�T�w5�����G�5��T���Ξ?���ݮ��n�9�"�}��[̑r�+c2�4��t������R�ǽUi)��&����?.�q+}����p��/l�LA��]��F��u�_k^��U�B��a��\�G{�xw���l�}�{���ZFj>j�VH�W8��P?�F������o���k9�Npg;+�ʉ�&o�Y~N�]pn|i���*�}���Q7/u����s���| �B���.�Y掏5����x55���_�x�� S|G܅ʶ�R14�ߣ�'�ܸ��۽��n��'�_����:�$��5u�(@H-7�OQϤ���[�z�7��GR/�80ʿ����qp�?ӈ;�g�����rz�P�ޖ����y2�K{�oVo]&������s��o�w�YQ�bԥhG�K���K1�܏'��s����^�-�"�4�.^�~̫}��Rw�u� �T =����b����|w�1�򫌻��[�:�)l�ޤ7^�.�����
曮:.֭m�g�5m(�� 1�Q��ۜ:�6�>#{}�n�I=ob/��/�'��Jo@SFn�-���5��Z�ٺ��J�K���6����>�ﻛ%�E�,�(��fA����Z��˨����v��J����MMmE�X]���˶{��+�e,�g���%Zl��Y�4�N�G����x_&ۗ��vU��q���y%_ga�����\��c��lO�w��Fk������k�E�?!��-�l��?���4Fybsrsrbcu�Ȉ70�Z3��]�r�5�������N�Q��\�<���V���ȵc�����۽�+��<��¡�ӦϙY<��F�O�F�[j�Q�.aC����w�����]��0F���l��X˕����������T�2�O ����Z�X�]�8�e�	������S��Y�0o�f�5~���U��ѻ�]�h�'Bi��z���N�N]~�M '�|ҼZZ�Σ��#�Tߡ[�s�(Y�n��7�X����yoB���������-��B��}�%���>V�\����$eki�h�V�s�me2B��ll�@���˅+pÆI�ip(��ϼ�����M7;�:��\�4)U�:xŊ7���Ds�m'^>ꢼo�b�iv|_�F��kE>NQ�4̾JܪܵIjj���Ճ��w�H�50�yom}��ysH慫�hIAK���緘ʂ�@�?��E����w57>��Ыv�E��(J�����%Gf�c_W�v��M�Ɲ��;�j��X�λ%*86�;9~�f1X�#��y�)]U��KnpI�R�|��� }�1�J��9u"�3��L�Ě��jl��$j
�����8�w�����8�G����MV�g'j	���r���&J��'&�h �o�J*jō��PK   �x�V]�!��	 &	 /   images/98931e0d-18f3-449f-8fca-8d5f6b2df0a7.png -@ҿ�PNG

   IHDR  �  
   m�y    IDATx���ٯ}[v��cι�ݜs~ݽ��U.W�U�I0q<�BB��_@�ސ�0!!�Ȁ�O�Kx �
&cP�8v��n��~���Zk6������ܺ.+�����9{�f�ٌ����'������n�Y��J��8"�� �ϥAD0��96�g�5�CS�)� �B��I���|=Nq��������eJ)���ExԦϷ�4L�Rw��un��p�ֶ��k����ᚇO���� �n��ϟ�{������נ?��&���#tz����ܟ�O���~͇�
m�МhT���������q��8�9�[6`_y�旿����K$���S��R�X�>�ι:����¡/�g����>NHh�Ϟp��������>�Z���n�0F������[o}	�z�,��V����X�����<�M�Q�BɅP���;��ۿ���a*D�Ւ����_�k�����D���%Թ��ȹ���iN���G�2M��	�_�w��������O^���f����~��_�*��_�m�]Թ/����E-���������_糏>��O^��i��8e�Ւ_�/�K��� N��ϱ?��<8��y�Ա+�����?�w�<f�q"��^]�ą�����S�տ�7H�)@�?���d�c�p�ه����_��|�=E:5..����5�޿��o�;��qn��)�������D��s�o��o�;����A�BX:6w�a�E����_�����i����L���b?��B>��9;	�[]{���A��m�S�������?<
�����������O������Z��t4*�?̌.% ��s *UE������z�@L��3i�u�c�B��;T�T��͌#)�c{���L���ʱ��qϬi>��?���99_�y����)?�w�������!����{>��g[�Lwj��?������?|Ϣy�����M2�/�Ə�nu�咏��,q��E�C~�{ﾇ�|�X��3OΙq��Q0�@��.��D�@+�8V"�@�>�����	��9M.��ՒO.�ay<���������'��,It�����G�{u ����{�s�������\1��/z>��w����'Jp,��i`������3:��NY6-ӓs�s�<ߝs����"u��s�up�:np���@۶�}�j�`T!�à�u��p��)H��V ���WG��f0�Sf@O)1���l4MC���^e*�C����ß��ID��9{q�`?l��-N<�E�>��1M�z��NA.�?�!M9��!�u4MChZL;�T'v�{�jޜ	!pp����Os�r�ZB�kb���GD�l6��s�9gb�x������9��0:V��틁������?+�����s뿎?��oց�{Δ&\��JA�Be�L�y23T�8o͌\
^;�i��'��_��Wy���g�8 iē�ƣ�kXh�1Bqe�Ł<l��8��Q��� j��?�Rʣ�v0&980���@�͑�9��hm��=��p��y����Ę�J3D/�b���Ū��*9g�e�v��H��p���V(f�\�C7��ѓ,YA�h�R@E(�g�3�!��Ӻ6f�n$H�֔���ɑ>�X�K�BZ<�G��6gid�O�ֱq+���Li=�������&�6��)og�%�5�!l�R����,JD΃���52��5{iq��#��	�)�:_ssǓ�W���ػ�\"9O�����L-e}J�u�b�#t�(9�_�l��MN�y�Z�:�<}�������>O?��I$Wh��5�+<�"p�k���u�U�6-�TGl��m=�WW,^}���a����䄮�Q��p;�����iK��	�y�E���J�{��A� �.`.��EB���eh�;�1�����͆��Z����(�ϟ���߽{�*N4>П�V�ZN��|��4!u=I}~J	�/�WGN����m���+޽���Ś��^,{l0���L�z������4lp��( %��� �� ���Q�^�%M8Q���KfѶ�|�]L;Yp�4L�kJ��I�[+䜑�%�@����՗�ia¡fx�F�f�*d��V�BbX�d2v��������k��;?&5��lw�_b�5"��J�ju�T�R�dC�R�s�<�xJe��)���J��A�)�!���{����e�Y^N.�Y��D ����_u�w������ ��*�`5�
i���9X�3���z��3�6C��6=���v��9ЬN�1@���6�{������D��p���,��_���R�88)P�ζ*R
��{Oc�(���eČb��8y�^�q����)󑢂D�������xþ�&%GҰ'OC�#����3yHÞ2�H�'�͏�<>灙(���H��!����ȎK S�_�����~�0�ȥ^�6;Ffz�����Rp��?��Da�6��h���LUi��64�l�<�(�.��u��#��<�8L�
�Z�Q�N�%=S�G� �t������c�JD��-��,�5���J�~0
s=~��M#���>y�E	�)"���EC(lF?G� ��B��%� Jh�㖋�s����%˳s�O����m�oZ�6�z!%C$$��8��q�R����q,�3�(cJ)�Zx���15��"x�a�n�D���iX�{|�Rv�q�1��r�e�G �T �q�F��Ǒ������q��(B�z����BO��Y�YOgK�B!��{|��o�w���2�W���$���"%Sr�sCE���8�h�5y�©g�Lm�+kRtd'����!���Hiq(��V#��=�J�IΎ�4R�2ىe뛆M�e���?�a(����P���k������>����(�;Z2L�lVYw����v^�s�B���V�g�=%f���i��ܰ�J6�У.��ړ�����o�SI�I�o��
i�����o=M�Tv,&$l�g�
�H]��OLˀ]^�b)|���>e�V�gn>����7��/�\؞�M�2��0�ɶ�Sh��֪s�&�tX��BSY������9�A}��Me*L��{���W�*�{����u�����'��u	-�=��N��-���
A�]a"P�PC����;���h���i�=9�=�ח�d�⑒\ype=ʃ���))f��Tɬ[��^t`"�a��2R��;Ԗ��-)*�x�,uU��Q�xw�a�'��b*Uw�E���q�ѿ��#Y�T�Xp)�c��#�<�C�������c3\��-q�æ=��7�Q���q�>G�'�'���H͉kzL��i&})�9��t�s�&*EjD T���n����@�׾��E��� ��X�Tf����M+���=)H*�PꠗRj?R��͞���c	�$#�4���RA�ҌMӠi�j���L��q@��z��R$�B��K�"����������T<؄S��r�i ��H�Վ,U�Qr�l�$gR��W��-�~��|(�GWk`q��#��4��SBJa��A�a��@�7�#��Z١8NL��J]H�F̔�����S���)�nO�7D���/B�����I�
*F�+jR�nQ#G'�O[bP2��y��i�$	܇�Y�%K�8[=A܎m��}��2�TC��`�w\ǹU��3ͬ��AQJ�`��&�("�3"e�H���z��%�W��'�GN��u�RX�)�����ˈfJRd(D˷�!��
r�HRS}iJ��S40LJzñx�-��r7��c����mb����G�2F:����H�9�����ȩ�HD1L4D�$w���A�'��jV����2�bÖ!��#/�������]Φ-�tS�\*���2V���5�H> }.5���I���_.�B�{��q�g%QTx�8g��m�4�𼅳�>au�)�*�\1�:�:���Uj�f��8���!�
G�o6��c�qN�Nr��H3�tH_�������LNɘ������t쬂�Y�����U�E�,�90
Ց�5s��1�zLk�pu�+i��x�xWSw�M��^������ih���	�Q��H�����]S���
�- �B��_G}X���9��̱5��ʜ�,��� �iCjxW�Q�9<��ӄMK�9�h͎��)�gs�@�Fˊց-��`OΔ)b�c]@��ޮq.� S�)1"�D�{���i�aӈ�T�-J��˃$��r,��懜��+�)3����I,x��T�C����@�S¢cS�,H)�q{�辔2{��}��!M����*F2�N� )��i�F&��1�k&[��(�X&皟wyä���ɒ*SfJ��Rzd�50�K���K6�;L��������2m���Wtc�"��by�D��ip��]��x�A,F2fM�NqM�*��٧�ݰ�����D[�Uh)y"O{�Ғ���c�f+�s�M���H�{(�)��c�IC<wi8�s�9�c��8��5ۻ{�8c!�X�i�;!�H,5��
3���ց�N�J*JA��Cihr���!wlr��.r#�ɱ����������y������2����Y�Y��a��i�@��>�ɠ(W�@5�#�}�b)�7k�YaW �Ґ�m�+���B��7��>r&욑\W�����ë��#ku|�S��h2��v�rOםs��5�x���ed�:��)�A�Ú����"�R��M��g��
 �Y"�LJ�7D�
�S*t�y�l�{��Ȣ#��0l��e`c}�w8�"~��*��H���3Й�us��#�L,�g3	��[�goٍ��zh�g7-(���j�8��H+�q_N�̟ո�vXל�ȇb9�áu��:�@�����vH���FLs��@���ˊ=��]�'ل���������jKƩK�N�%WG�L��R���1IŎ��C���?\{��t��Q[SI�YC2eQ��:�mZ\�&��g�{T�Z�oq.�B�oZ��pQ�O�"�!~���@�5�m�|h��	�=:e�i�0E!ˈ�
T������l�����#�s��^�V4DD�\�XAb���I!{,x�GHӂ��-i��b��ǩ cfX�J�'""�9_;�j�U�'�>�1f��IumP�-��=�U�LR�?O�����Qn�$�:.���r,Vʿ�VY�jl���w8[�k�9M G�U���x�@K��9���T�\bҚ��
�(	�~�m�nɥ�٢�BpӜ+w�;����Hβ_3�ݱ�r.���9��}�ܩgg���pm���RY �"E��
�2��clbh�H3UUT����_�\a��xJq=�a˔�6e��{�i��	;?ct-��(����1/i
S�(M��-1�A]��J�25kr2T�1�K�:z9#��G��4���HQ%)D1R��@��t�-Z6%J'��H�| 9�]��s!,:.�>�iJLW��{̈́n��k��&�{�&���kmp�XR����!��W'd,��N��s�S戻˽C���s��dX�T�y��=>�X�l
c��ə�m%���M(
U��Jc��v��;�LFJ�X"��&��p�%�ἱ����5GɁE�bf��#�)2�¹_��0����/
�֥=Zǔ*;�6��f�K8Ql��v풮�r!N��r��6��4�F�w�����#�B��$���R�����(�PM��`��X/.����
�4�L[��E�X�<C�H�-gmGp=wS��XU,�YEfQje/�����~�η���W�G )��Xelʜn�ѓ�UW�M�� :���S9�{/n�A��I�tݜ&8��L�FJL@!t�����=)��)d���ɜ�� �N�T)�l'[�2^R�,���مS���Ӥ��Qf�%"tW�>T������6^"��%<���:MCj���aNI��-�b�����?�2O.^i�ęO�ua�����c����|3S�T���|�.���Ε
+ӄO�j@�Qy�\��<!9R��Y����e3�9g��x��K)�9B)s�c�[������u����p��	�yp=_'�)��ɇ��G@b6{jV��X!e�Rԉ��]��l�13��1��7S���69>���L1�����yr�Rtvp��x�K��{>ʙB&�F
�t�<����~�����)%V����,�q]����-g�'�3.6�!�%���ŞL��s�~�-��mj,Զ�GTH�	����3�R:�`�5\o�1��4��A��%|�x�u��&%4E\�jD`�Ü�ep�гmF����[�#R�2��MN�T��햱�����G�����%.���R"�#)	ΠX�@h��dQ�O�W� !���
��pa���Z����{ٳ�+�
�0�<��-"Ɇ�os��
y�h+�Bֆ�F��A����,�5n�8�&l���W,:�E�Y/zV+�4������w������5js��Y��@A07ӛ�j�W2�`�%��͟�v�w~�)m����XvkĿA����]��Ʉ�H�Wla:��7���:(#���j�r�����Ĳ�~�a��=c6�Ĳ�9��!����\��*HR2F<F�N.&�Ug/�RR��􏑒aΐ���R��e\3"��#������$�ٍJ��D�]��r�V ��x�;�Ԭ��p��!&�T�AM]�uW
�@9��T�j��PQBM��q_EEP@%��dTb��0��S��oʕ�*��ʂk�1h�1���j�c�U�>~R
�N����.Tvufzf�D	�+U^5���!vۿ=���j�Y������9��ʜ�.TQ�F��kEP.��X�c����-zJ���8m�\�Bu���ӎ�n�G��VՅs�H��<�p^]��a��%F�&�S�[
 u5wR����RE/�P�S=G�6'0�� �cn����6;	:G��� 3��!G�ёN���R;�?]'��?sz@}�J�<���Rr�i!;R���]vL��)A�TwI�Ql�mǮ^_'u�P�.-�U�(K��'�)�u����ߎ|:DJ������h),.����YO0�{J�t�������w?�#�@w3�kx��W��e���̤BRx�������u�$�u5o��p��(X)����~�v��L;J�4��6p�3�������ky��9s��.H49b@����]3u=w��}�f�#愪���D����L�pn+��1�&�o���*/S�zm
�͊7�L�E�i���#q�!�4���֌Ϧ�&+��Iꘆ�S�X���=gz�4
�̀�H\GB46�;R ����9��3:��IB?)�ThJ2e�Kųw�-�4m�O�"�zG[de(BX\��}�e��!�Ϊ�#,p�����&9�(|i�b���pZ�5p�����g���͑���H��g�3d�m��z��C�s��H�asw��g_�֯sռK�1�t-��E�2Ӭ`��b��Ȅ��[�d�)�bx��GD�Z��3Fi�Ii��uӲ�n�c��@4ϵ�r�eM�0���h�!U�����<�E(�c��y(5}'����i϶i(�D���K�빿����&E��kLMëAXJf�Z�n|�3sF���f���	��x{ F;����t�������pW;U�a)���0��0�ڮb	��p������*!h���DMs*��	,S����Q5��S�&w�g��D��1M1󢘝lvv=E�1�ef�~ Q�c1�!�~~����ˉ%@+5�K�;�1sQUא=��s��#4��sIh]F:ǐa�������c>~�熕r�4�b=�_�r�?k}�}�r(i)FN�]�SʄZ���ܼ)N��9մR�3��97ԟ�rf`��=8XG:h��c��q�[�L�j������g
��M����:s~��/��ةj�� �A��r|o�S5-13Ԝ���w�P��Ww�;ϔ���}/W=Y�M�T��1aL����yk\�%3�����%��L��O��KL�]�4�%�2UJy�ś�K\εL�<w�;�c+��n��Qʈ�P�
�nx9N�����W�2����    IDAT�)��q��*��G�D��!k�uB�	#�_�^��L�On�� ]��.����u�`e����$\�&>���h2�&���<ҩgMܓs�+�L�[��:q�>��K�9{)ܥ�o��2��M捅���V�Gae¢q$`?�:{��*���޳c��K�zC&v�g�L|�_q�lY��+_�;O�Wжl�����pyǓޱǅ��ղ�L���8>k:6ŸN�gS�6g$L�f�a�O���Q\�\2���j���H���
Ʉ���I>�^�5kw�[rE"ј�[&dΟ��_eS
W�x�`SJ�'�2R������鲰����]�I�ݾ�ɂSp�s^����j��by΢�ƏF7�r2H�EYB��tY[='�����n@r�c��Q�=6fB߰-�q�-�����o?�[,�(/�%�B��g�a�\�82N�F2a޿!R()��X1�LR%�sG���	�����oo�M�=�_2MB����ptl���ϑ'=qJ�fᙟ e`�I�;A}��͌6=�g��k� 6Y5p"�7�qG*; Z�D_�C,C)����h��L�\� �\�7*4V��u������PY�C�a��������Nf�Z�y�U���dRg�攩*���jv�����Df|��Q���lZXu��R��pm���,�����^�c�
(�u]���æ-;K�Y�?�p����*H�us'�\1�BN����R�P�f��r��+�lϹ�a�0�f��ۀ,��tRVd�|��+��v���p<�9��p �CT<���I�q����9&��P˪j�8�����y"豝��;��B�H|���ǩX�(�R��\�y�
3�\�� igE���+�|?a��Ɛ�g������;��~����K��`7�1�l��4���o��?�{������Hd��ifD�kwt,-��t�д���o2���C�X.�4m�k׻[6iK2�6��g�#��9_y�	Mp\]]r���]�nJ�)�	��,`x��:�eG��Ojޔ��%h�0lHe�\[��;�6w,�\�	|���|zY���&��Y�F�f��Ò��vSĹ��{Rّ���L��[��7�|�1M�y�1�����
}
�Z�n���g���4����V_��#i7R�5��5����W�|��p�����H��z^�#�@J����zu����bMC@]�^v�Y�,v?���G�-w�y�B�|mu�WC��%_�k�.,x��||}�g��^=��~�/�L'���i��e�\��f,�����Lnb��[������;�g�x7]�rT��*o�-n��L�ܼ�������y��CSFbU��s��ٿ��m���mu�qd���]\��qB�c���{>��y���7�|���C�_�ka���X.���Ƈ�u��������n�%O#nV_�q13���z]X�S�e��eЉaJ�����Վa��������g%ƹF�Y��ı3aߴ���v��BqE�)ML6bR0�ȟ�x�<?_�v��#��}J�N<y��}���VI���Ο�|y��}�k��|�`��D�L7W-7���;;U v6��ϟ�Z�r��nf{1���hqvT��ys���x�ڣ�%"�Ӊ����R��FƵ��������,���`w��i�jy�s����{�Ĝ)�!O��y�(S�spQ����%�P��(9%�k���F�<Pw��2Fe�x�8T��Y����$?�����x��i���pQZv��0��B.�r�w�R`!��D(�㞈&3�},�8���9������vl��	(kDz.��!3U%@���IP�?M�?8�_��W}�ó���j���͞X�Ϸ��{9N��a�h���|����t�4��F��X�Z���+�#3�\��s����z�������+,���l�;��x"��v�|�����[G�e��HD\�x�'��11i���z�V+.oF�8�Z-�+�С>�4�؟1F,dB�T2Ӹ������ʿ�?�?�!����17L���+�N�j>�BT+8�Y�K��E�����=9����VOx��5�y�C>��CBhx�K_b���L�[�#S���+�_��W������}�w#c�DfGl��Y�g�������4�s�������l�`s�g�߲Xtd��� M��dhi����7^���ow|0\m6진��VF�RKm���6��Y�Um�Sd��!��id3m�03v�@*�����Q��|I�n�Y_A�4�}͖ͫM1RӀkqA�nDfcEA�⻖,5�C�l�W$;�EOӵ�zu�vP����Kv��Yvąp�xB��,��;޿��2�"dW����s��W�M�#m�3;V����~u���]̌���jÇ�7���=����C�~?�x����n����l&&�;�S$Fb�5�ͼF������H��_ֲ.���\�ݲ�ݰ]�a&\��WCC/���1.n�wyy7p3D�$PG)��D�BˮR���i/֨w�]K�Z���~�	V`��>�b{w�X�Onw<])y��m[���ŉVg[���cN�`w��';��S�urrP�NL�ц��Ս���ˬHw���R���?��pN�6�D)��>���f��P��d)2ofS˫W}�L���Z˟sƒ�]���:1�"m��;b)�o6<�e��蜮�X.s��gr�aWO���f/���'�S͒��.HF��Zi�G8B!K���z(���b���bN�5*`c�z9ֈ(��J��V'����[(�Ò�#~�睢�Z�2�<1���� ��gG���G}�Q'���E�8M��5���Ŭ���Zt��Z�����;�`]8��I�2�p�뙾��
s�dV��πł�H��j��_�X�/q��_棗�X��6��l�����G?�17��.^�6a����Y�dI�B���;�j�������+���隔���(f�)�*4�'4Ӵ�~M�x�o~�!%~���}��g/�nk�9�'�T��T-W�l�Z�@����X-�<~�j������8;[�|����[6������?G���?�>�����a�!����͗�UU�\pt�#��J�JA��K�sL�O�W�SJ���QI���@p���?��������~�ۼ��p�۳-0��K�h�N�ֲ'U�q���n�j�̢	��/�q����`���e�_�H��hp������q$�W��_�2�O�|��w����U)�!P�-�z�jJ�iD����е<��ct��m_��O^]b��.Ϙ6;�\AۖwQ��g|�/��k����?���;S��PZ<u�,U�LPM��:�����b�fL#Y@�c3�2H�s��=FG�	q�rߴ��cݚKu���w�H�CաX5�N�PiԶ����m/��!�\���Eц���iV+\�f����8	ow-�o�Zŀ��\i�G7�܏#�@hjj�D��P#h�{�j%a�Ⱦc��_f�����Ħ[�|<f�����e2�z���#,c����,NT����!Ӝ1�ǁЌ"��A_t ��ח#x5����Y�C�k��sm����2�^���T)���P�%�Gfת�O���-�{$<�(�o�@{�Ô)�,/���I���T���5�b�64�rb5,+V�.�"B7�	(�� ����0�?��&�Y��Dg�Zͻ�o�C�RS9Z%W�/u#6���<8�i����A�W�� �O�w�G�i�h��_�pV�m^,��+�IUy�j�t���=�4?T�;	%~�^v�������>����|K�F돢o=h����V�㖴'�*G�8�/َO�� >Pa<l�\b��#�L<%à�ܮ��������k>��C����;\�ܰ
Kv:�I���:��(���O�i�q��B��«��lE�{.��q����a����;������i����7Y_<�����֏���/�߽�68�F>�Qp�2��5����׾F���xƛ_~��?���Պ���G�������x��^��j�|�=~��w�-��)��[Ɣ��t��1J�1G�Ο1l7�������[����W����p�ȢܺD�;�Ӏw�l�X��چ���������t�i��8�r�R `h|ӠZ�Ip��o�,%����g<{v��Y�ۜ�V+�67�)�G�)�}�H]��O�&.�s�g��_"��-�8FR�������qJ,���_�a�X�|u
���W+^�zE�-�E��J�[�e`'�8V��^���|��+>��ڎ����y�\jy��RU�J�Z�EeUV�m��O�-ȥ����'�XS��t�#�����I���������}��������!�4��	�k)N0M�?k���Yv��}N���'n��)� e�hɩ����%���v) 	� ���0�;3;��n<�?�{�{���T�SS���Nx���>!�ۆ�b1A�%uSBc���l^Pu[Qv-I��{O��J�|�:�|����I�X�zΓ�WT�$� �l��6�s��I���� �����9��`�d��ޞ#�(�-�i�W��l*�"�	H�EI����!��3҅�k/G|ގ��o��;N1b*����"mm�� �|�CD4Ds��8ki��Zӳk+�ᑺ�����	���L%�������R�-�ơ�:��m	�3�rO�������{�"�
g��#<�^'(I��r�8B�@�M�<
)b��
�u�h��5��xgB��S����\c�7R�:������6�C��f}�l���|_�է����T0&������^?Ɵ�C��1�|<��H��UT�}�{Xl��7x+Q�Km��\��$q��fh�p}8� *����f4�9��D�8~���@����4f��C����&>���d��-���=��O?���l����g�����͚mSK\(���(�l�l6CX��j�$�(
�y�]�ɟ�1W�5�y��w>`6�a]�q�/@�G�d��Qnj>��N<Bشh����g��/t0�T����QKE۵h�麆4�����i����GS[T�����?��@(�D�-;2�PZqv��=Y�"\ƽ�]�p�_�l,��g 
*OYn��9�ł��ɧ9��.�vK"G'��e>�SWN_='�@c)�E�eO�y�ݻp^�op2%O,릡u/$z(A�vl -i�ɋ�6�f3>|H�VEZr|'�]��b:����quv��`��C�3��W;��9�����	tM����S��f*��V�9�/YS��tXہ�d��������W���w��n:�>x����/��eY�|��WOp���ŁUL� Wo="	�;cmh3���{	�;��!�d���'Ֆ<S��!,�����='�򜮭� XW���L�G���k�C�i^��	M�O��Y���iQp�< ���1˦��%��.�����A��D�,�qƓ8ϋ6ᢙ�g
l�;�V%���=��%x}h�3���cڶf6��u p���]�)�w�T�@�4	ev�q(k���H(RZ�z`��ľH���Ԃ�/�P�u奊��X��l�2�p��dEDo�Z�a{���o����^�w8l0~���2�����u�d�)�ڕ�U�d� MvuM�r*�Ҩb
*�4W��xH�ڶ���|���hۖ��1S)�	���)P����J.��~O�1M־��:��	
��ӓ��#���s�cݟ�}+T
�a�ayp�"��-*������y�ȷ����̝_+_�_�C>��b��>-�[|X4�
2Z_�s��%F�{���>"�l\�ױ{�fT��?��V���:�7���u���{_��n���� �U�7�@	�tL�cc[���4a׬y}��/�>�C�"Is���I� �R�Ԥir�Z�uOg-iVp��}�i�|1%��U,�4M999a�m0]K��䓂�g�y�>'M5�Y���f�K桜S��#cF���O�f�u�j����1�[���X��U��'L.^��	Bv�-�^���?���g<�xŽ��`Rx^�zA�uHB6o|�怴H���b�r6'U���S�=�Ǐ�c�������ﲘ2?8d��	��+�ph�1��v���D�Ȕ$��sh�x����2pUkz6/�����9���?��ѵU0Ȗ=x��٧���������OxCSm�w��,4m�� ���i����KZ�Q�`8���dRTUE��p||L]�Ȳ�;w���C+x����^�(�Ie�i;���y��8��@J�|v�f��n[����
���F�N$���G�|�{�������3��=���he9}�r}��-�`$�<�V����彷�fw���l��U��^��ң�Г� ��t���L�����?�ږ4�`���e�����C����Sv����ˣ��η�Y���sLՑ,�Ts�=���ִ� �'I�p}�h�C
K��,�s&y���=l۲Z�X̹l��vK�k��&��1�%Rv�?��#LSr�ې(�Lt���{nOP6=9�^��!�!�/U 
d(���� 5z����>�A)z��y�	^�N�R����&Li��
�e苹���YJUUH�ɳV)��Q�R[�FO���wx�����a�+i�3)ft"Ȟ�nX������뚺�9T5g_>����!O/9R�B�$��ڄ���5��t-=8/{��h�8:�P�b��v �G\B�>]�]9�A�����*���ZD�X�~�k�����H��A�~`#��]W��{e"	q1��#��H&*�x��C�k
6>�p�ލ�i�&}��h���W}�h�J>\�+�D������P�)�;?��*\�?���G/���4Nk��©����C����dΫ�j[���L�X/i�Vo�����H��%$�/��]@Cg9�|A�ͨ�-y��������)�{d���C& U(�L��<��������ìH���ł4Mq�!�$�3�$a�d2�:�&!�&�EN6ɐ6E�P6-Ƈv�����6��n6��v�g>Iu@�v߈��_,Y����6�Ҿ9���`�����'��&MC�$�	D�鄶h�"L���O�[�M�?�0���	�+���>m�BW[cZ:�2��x�[�!%L��ɝ{d:�}�y�"�#��ڃ��-���S�~��Slۑ'�Ty�?z�L���a�t�bڀ>N�kU]sUW�����]6��r���Ϩ���|��K�#�RR]�y�V�Ֆ�N_���C(8I�݆�5�B	��rJ:t�W�I�1��'�dx��#�|?���F��4q��_�G�L&9Z&�"�k���5/����ՆDH�i)�kL]j�i��A�8�>��f(����w��w���̖3�'���[l�g��x��-]��F��r��P=x��dN�NI��W��ݮ�u�<Z~�NH��$�@�*C״�;ǴuM�u,��"LC�����C�ʩ�k::mq�bv��T�
_]�/^!���D����B_���5�{$�o��C�mpC����@��zY��U�H-�Dm��do`D>��`��5�u��ù=N�h*�]�P�De�$�q<oŃ�y�?�уw9�s���{�ON�Ӝ]�ruuEYU��e�YV�-�U贘�9������\s��]��P}����/�öb�{�O��'���I�7}��`�<3���ÚP�J,��|@{�o��������Q�n��Jv����׽����p��=c�����������i��2��3	/�蘣�9����_=��)��;�r��� �>&��8����DP�5/�/��}�z�S5��(��	3�C"-��KD�H'�ͨ��i�ٶ�f��w�ń�	�T(��6������"�3&�	�����i>!�6mMY�$	t�%�2�ے��fEhT1�Ni:A�ِ�х�Ϭ�a\ [ҢAx��fm��G-&�����T�&��3$Yʝ��8���ͮd�Z�u-�̱Vr8YR]lP��0/�.qۙ>��W� d`�JҔtRP�tU���%�������# .//�u��ߔ�錺�R��y�� �%I�v��uM���\m�h��&���M��K��-D�#����)i�Y,�x]��7LS�d:�ZK�۠�&���;'خa�l�v �@s��A�mUSi)��    IDAT����	�;ʦ��f迀V�:�:^I�~�������k��9��b6�ryy��lRк�@�͋/x��y6��0:	5�^�|��sf�@K�����sx�$K��	�9��;��]�e�I&�M�b����]g�+G�=O>��O>��`>��t-uW3���t5N8�D�UPB!ʖ�E������|�מ��#����d�sy>��� ���ѩ�KM��\o��o>d�N�X���pvuI!Z�0t`j��$Y�Jl�iMCY>!�s��	:My��x��������������$����j���R������͊;M�ۉ�Ӯq���Bg� ��k���O�����%�Mc��#�"V(�k-]��xk�#Zj�*p�ۇ��k��� �>4�F�J,E6a�m�U��;�������$w�q�{�O'L�S���/^�����/�mZ��sp��*C�!!��i��T��Ӕ�2���]f�哯����z7���P���p}�����t=��C���)�GE���_����0G�H����Bn�D&%R��QȆ�S~�Bˑ�s���@�BJdC`�J'cN�wأ���zo���t�=��`e`u�^ỰhT*Z����~i��x�+G����}�G�
X�O��uX�1'�F��W�2x"�h9X���ۛ�Bt4���95x��{��Q�����Z��H��5�z�;C���n�8
��x�3$�;FIO��J�i�{'C�VY�x��!�^�)H�b����PT�3��)�kY���Ԍ��D�V\���a}%C}��o�#I2v��o�hk-��=�XR+v��bF^TMK�$8�pԠ�u��&�]��ؕ+��lw%��"f�!�B�̦iȲg<���F�r�����I�Ѹ���C�d�:��M����3��Ϲ\W���6h��I��|��y�=.�}��t�]����Ӡ�
	*Ѥ>�XLX/�n�x%�YSd`�,ϸ�����#.��w3�\]]�$�8$�4�b���,�6`+�$�{*X��=(f���霮�m��,'��u��k�4����GW?G���,�P�J�$I���ٞo����D��Exo�A�T-�+������{�c�Za(H��1�t+Φ$B�f%xO]�zC.���2�´�iȵ��㲡�LP8�$˂+&9<`6]���;�ܽCZ,����#�MK.��∫��w�Sp���9+6|�[�mX��WH��
L��@)�$/��J�?|����8gX]�sr�?}�m9>)8�+2�`��=^Xr������Hu�Ʈ�N�YF�k&=���C�A���7䙿|��|k�]�N��� DY��(Wc�҅C��wv /%I�t�h$6�T�$�)t�ٵ[:�9u]1�Mظ���ۤ|��w����>��d1g.eY��/~�W_}��O�Q�%������|�H�~)��6������_J��dJ��ȴ���'��b�-��H�E����ȴ@���!�~�E��6.̍st��iI�Rh�2,��+��I�p��u􃻼��BG*:���Y��u����q�x9*'�Xr1Zo�|�Ml���{7�V��T�:���_Y��Wz�N�ka��5��r[Xh����U�2���׾w[T">��A�ct�m߹�}7@Vs�i�l͖ �� �"���J%T=��ZKS6���%uc����G4B�R)�����5��4O(�-^i�|2G+�v�e�Z��c��!�*�B}<.Q��0u �Zk��%��r�6k��2)
D-PiB�'t�Ex��)��4ϰF�fI�oj���W�hh���d���!i�ruuE�6ܽ{)�_���J����)��j-X�6쪚�d�v�BJM�u�����AJ�r����P6�mK�u�Z���,��J�*�	y�4�AK�x�~�L��	IֲݔT�s������a�^���@k=��g��t����n�֚gO�P7;<x�h� �H�u���@���VR6P\[߷��o�C��4��k^�z���n��H�ВX	2�;�T):-pe肨�C�.����\�\���{9�)��wam�`-���䰶�jvxip6�/9�^[�c%5Do��q�Q�K�I(�������3�D�f9���iC�ll	�e	McpƆ��I
B`[�i�N�}N~<}�r|�O>���f����-l?���Zf�%u��ؚ<�(/1�B�9�i��������`��?��&�{�˃C������׿�5����	RK�BIK���$:�������=����CZ/��r�z�e�Zqq����9m����G?���S֧gd�AIE��$��4��s��u*z���8��\O��:l���m1f/�Ǉ�80�ư|T���m,Ay����a�W?VB��\�{��D}ӤŅ=^Cn�o2�������Д����$���co������ߴ(��uK���h�?"TaS=�m�)�G�zr�2ѨD�mm5B'��;�|��gϞS�Y>^a^�"�c�eY���b2���
�rE��\�רD�t5W�,�����rM�d��Ek���p��sE>�<��b<��Q*l�J��a�XPU%��:x�^����M����Y�פɔ]Y�ٟw<�qB���d2!I�.�R�޽�5��,9<<FAӒ�J�ФIhN�/ٖ-:ͨ����@�yC���5|QɎ��9G�e,3��K��Ѷ-�X�]I>-�:�
^�:��tE�v���k!�o�	�ʾ�D|�i#4*����{��}�V���K����,s�7��8���;�(�KL�c��S:+��ӷ]o�^8�ł4I(7k�INgj� U�s���%�.4�ބ(e�^����a�0���@�v�r�~VeE��Ӷ�$�F��|��J�VgH	��2+�ɗ�)ʛ����̒R����������$I�-�Ȳ�������j��_!bU;� UB���5�ٜ�4G��̓r�b�A�EoC��9�!�nzHV�v����:�lɮ,1�R�9Meh[��3�(6������Dw�����#U	��������/^�Ѷ-y^����<|�6���c�^��'���÷��m����)����)B]_R�5w�~�ښ�披�3��N_<�$G-��+6g����,��x�`}�"��+W��:>�'T����hq]�ao��@z�A��p�冹e#�K�b�W �9o����?bӻV���w>�������m��vV���<��J�К�Xg��~��R~cQ��oT��Ɵ�&~ |7�7m���k�|��[������ѩ7oo��g���J�a�F�ŇҔHH�+��tJ�=W�@�+<ִC���i�Ri�R�-u��Y�t������HtF1���l����/^rqqH��3ᮿIH�4��l��sǉϟ�)O�<���+�<��Ζ�l�8|��c�,G�z�C�j|��5�s}�^��$	J����׬½Um��	'''�����Z1�Nq��dZa]�'�{�j�C�c�%����?(��>�1��7��.��tm�凶�]ױX,��a(���mI�*����ϸ����Ɖ)4m�޺R�u�Q��&���TeGW��͖�bA��Hf�yN�*�`:>{�5�MKQ�L4ee��vH���~�애��<�����ښ4M�s爦����8�X.q̺�Ͽ�j�B�s�w���y����PJ�[�M��g��{��-\.�LӜ1�:�I�f����+���f?��4VTC�T)1�bܾ�$G�iO��0G�R���f�������yG��n[q�ڠtJӵX�Wk�%�`:��Ť ъ���辩�E���1^[��J��E!��QZ��g�ɒP=���Sf?�!�I�w�=`}~ɿ���y��1Y�8�s���#��������l��2.OOy�?���{��Oz�iYoV�z���_~Ƌ/�K� P5k��$��|���;�y�}��w��:�z�%��Sj�~���i�K����LgC�\H�XbkL���F��}+�P�G ��aJ%���n��X�<���� �{��a!n��5��us!�����(����w}�߇�t`]�C�֑$����֒$�����`���`���oz���
�� ���?o[��H���a�po�g�{%��J�V/�J
ʺ��R<:b�xZ��I��,G)9xwQ�l�[:g�r�����9(�SR�X�w<}�����@���b�AH���֚��[�=�&rg���4a2�!t³��s~q�b���v��ū<}���uA���k���+����TTm۲��k��?>>��:~�˿e�Ysxx�Pppp���)����ڣ�N3�>k!�0b�pT����7o�c�۱Y��f�6%���$���e��&��K����ڐ
麖��0^W��?��YL[ �P��!w�a�4��X��=�3-���O�'�����_��%TuCey��4`��ƢX{Z�~���~�?��-�V�i����͊b:a�9G!8??��ӧ4�!����o�A���P�ؾW�^1�׃��tJ�c����$IC0��������E`�%�Y==�{Л��W�{�vlp�fiV DK'��m�n�cHӔ���������B�X��BZ3�
���IU��d�D[l�C��s��{�o���^��i�=���18F�us�{��_W��H���y2�n�����6˟���O~LcCc������_���xa�|�>:���~����(@(ʺ��\st�����n����|��ox��K��K6����
�-�m_�7-&�99b�\���?��'�{oQ�t>��4�<}B]�dҠ=h$�3��PڧY����>M�슰/I��!����,D��Hi�+�X���B��L��9����8�������X{N����?�s��b7�����t��,Kt��p���I�W4��K"��p��5����B)�Q(+$�|\7V������W���Y�{GP�} ��a�G���?�!�XZ!!Q(��}'��vKWWX��B�"����M*�$�1�d�u.Tmn6(��珹��������9��Xowl�6xQt=��g���8<Ǣ陯�в�碬��^Q�&'��Ϟ���SV�U�'�/������)I��ޔt]�tޏ��cAs�㴅�A8G�@�4H-C."�-.W\^^R�J?~�ג��N_������=ۘ��r���r�.�`�4M@�������*���Y޿���+�<�2�l��
���ׯI�9�P	ɵ0�s��q�p�N)�0�i�Z&�	ƴ�m��rNUU|���c�Q������|��K��!�m��)y6�n�ў�ݨ��t�ǚ������>M�����Mɝ;G(���ً��:=G��B�w��hO���8��3>�͈BY�Czc>����K�Ԝa:�����XoJZ#q^^��zsƀ�q�'�r������rN_<�5�ɬd;����|�ٗ����l�y�h�+��-i;ѡ��v5�u ���!b��H
�䳿�J2�n�!��i�b���O�9����/�5s�z�]>�����_��L(|���;�������er��	eݰޖdY��`�s�������o��7|���֒Ȍ�1x���%[W�T�`('I��W���3^~������wO��g�,��WO�2��Ȥ"���@��ߣ5iM�%��뛣��E�v�#5,{����[��q�pC������h�����M��)�h�TA��E鬠�#Kd<�4�88:�����Fts�����FA�}z��.Q����(��.Ⱦ)�p��x�{���g?t��i��ۓ0�s}pH�
�Q:��z��1�+��iB��:��8�sHc,����:�`�]n(�הe��AA��!<mW��� �����1{�7��9G��U�4�y���d�	�mM�R�9�]�/[��A��r:�ݘ�q�f�>*X��L�4��oۖ?��]��v��zM��0��ij�z��9JҬ�v-YV\{��8���`�D�U!eYrp��z��g?�mېjI�%X#�-ʦb[ux�A�-�s�ТaS��p��!� �B)eT<Q�V�$ih=��9O�<a��QS��wLK����mMәO�(���?���� ʚ�w�T�s���{t�as��nJ��p�<(��>~̫׫�i|h�26��#���8>^7�Vc4�����9=}��`���EH��_���+�^�lt*�+�qz,^w���6��!���,�K�;������d�zuI�%�W+>���Ӂ�K�6��C�*d�P��L��\
dۑ�X���:���`o��m�Λ�������D��\77uEW�O���E>�����O�9��c���;��o~��_|E���d���?����O�J���)/_�2_p��!˧����7����?c��ѵAB��(����H�����/m�:�,�P��ٓ����`����9|��L�3.�S̗�`�5�������7�ҍ"��2�7���A�}���z�H���=C[�azJ�'��Ľ�4��9~��C>�W"�ҵ6tI�iB[wԭ�[K!�7��a��с���m����D����^<Ͼ�Ի�E��i�k�9lp��H�{V�}���t0����
3��]��A@7>�I���xi�S��1���B�E�e<z�)9>>��$�������	Ϟ��9G�44ME���7��^Ր7�v�蜣m[�R,�,3�$�1����szq�)K�Nؖ;��X[S�%ǇGׄ'p�{�׉G4r�,�m�AQh�)��d�w4��j�u\�%��:QiG��M�d�h�=ݽ(uOOO���T�"G��_��%<m[3)1_�Z]�^wL���PW-Y:}C�h���jx��aLH�x���M�:(^C���Ǐy��9R�ʎb1�Ν>}��]MH�4(eH��g߼=?V�q�\wRN�&9��/�ׁ���;�L�K�%�[��q6��t�MoYa-��<q.i��B������>��l�Q7�pq^�?��U;������mF�M�?�����2�W�|�R
�<��Z���]my��5i�Q�QZ��L��鐲�Lf$Bb�ٶpZ{|Э��x��P����o� -l�Q 5����mNێˋ׼�,��_���_|�-2�D��?���ɏ�+�MC>-��z�'�~ʣGo���..^�˟������٬��ݔ�+��(�@n䤃��ˎIqL�T�U�5�2��Z�Ʋ^�9H
l)Ț!����޺��o��l����l��ė%��C���y�~���g_�'à��Mc�m�[�ֹѠƓ9�:�_����/�и��&����gJ�{B���'�Z�� f�4T���Q����{0�q$B�J˫'����s5�Ѩ��'9.
����!�C�@�r���o��"���$��u�q}�J��9I�R�~�q��s�������6��H��<��zsk-�N��3�Ɠ����(���dy���(hՄ��`6?�3�j(1>p�+��U��b���ۏ?C���!�%�o�"MS>�������>�R�-IR����`��*��l>��R��Tu�c�I�^��"���<I���&�IXo�v��6��G���,��c�Zs��	����f3ڦi��tb���Ѱe6�����劷>����g�X L������gϞ�g�ބ���z,Qy�OpTJ���!��Q�Ʉ�n9>>������/�2t�+�*�:%M<]`t	�.�Z����7��n�2��XĔFܛ���$�?�)'''|��G�e�NUU�W;>��	����r�P:�m�����X�GC">����]�v�P�v����/._����{wO�l>���j�h��D�&�΃�#(���C��[�����0e�%MS~�7�'(����ٜ�n���0��1v�s�T�ȡ1Bߋ���&^���i��ϴ��bz0�����m,]�0��Lg�ْ���૗��Z��j��:����J����;���t��d�i{�=:2�����M�&��6�~����C�ػѹz9��2���M�̩�N
i�ڢc���,�����QO�]~�F�˗kʋ�dAUV�7�~���-�i��2�ӿ�w���;<�w��������Ƨ���y1%�g�X�Q7�3}�Z"����'    IDAT�5uհ�O��MӔ�t>TedYƅ�QVS[S���l���9�i��O�����RlZt��IO�:�W����H��@xM-=��v£�:rCS���O�>$�F��C
>�V��wmBś���<��,؛yCF����+θq�go��6����"��6����w~E}Y������{��,-�7S�0���o��o�}��m����xR�SVkÎ��%	^@�6̲�<�N_pVK��+�T�hI]^w���K������<�͆�
��� �ggg}��&+r��a���4��0�^(�8<<��p>B-MS����8l0Tϟ?��t{��1����l���HDT�u]�eِk�׉ ���#2�{?({!IB�WWW|��G�5���i���Z����{�yo��5�"��N1�/�{��TU�j���}������H\�1j�6q~�e���U)%�x��p�������1���������#e��S7��=�ۼ���hL��>J#BAyn�k.//+�%�3�>��%i��]�f�(�M�!w3��g>�\�Z��4�����f�n�{�<8���7J<�H~Ƶ2�8/RJ��{@Um��S7�.4�r;϶ڲYW��_P�u��v��,�0HgCٱ�L�b�r� mh�u[Z�c��ߧ�ǟ�&����õ4���� }��.��s������?�}��OY.ζ�a��_��?���'�]�Fx�RͿ�?�W�K~���_|�_��_p���I>���j�eW��k���\{�{"tl�C�Ά4c��ߝs�_�RR�:�bۆ��=��9��|��jK��SvMKB�o�Ь-b�`������c �yݢ�mBƊ�^��$��J�nN��>�mo	k�?��؉}��������I��Fl��O���8<>����/ٽ>6����aD���K���Q ��׼1>��[7�M���Fc���<��I������n�$=�C{�R�7��zAWbL�N�s+A�Q�o9A����Z�d����WWW(�r����l�e��4�	X (e�U���d�r���?��ٶ-�_��I� ���jW�t�^�s�Eq��i��b^<F"�&*�(�gj> 䪪�ZK�����4�?�����gL�2Εg�!����Z��là�:������E��>X���N�Ьh��_�' T<{���o�o�����n�DLM3\�O�x��e�k7����M"��muR)�A����C)J�J�{����ơ��5���mȑ�/�͊�� ��ȪT�e�n0�@Ƹ������|�qzj�������
�H�4�զY��)BZ�z��V�MO��h;�����6�YƝ�	-)a,Bݼ���v|/���m�o:��8>�?$5��Լ�a@S_Iԏ�b���񺳼���8&����	������gXk�M�������_�'?�g|�����/�ӯ�pttD�����$@���j\?�RF��= �i�aM9�����u���U/c���t�}����Zq�B��5�}g ҲҲ��zC��~�)��D	����ȋ���>I��;�/o���������>Ї�����㚸}Q�`Y׊�NBd���uf�_Ӽ�R~�5fS�OB'��֜s��5,�pS����h��a��k�{E��[�9~��&�A���c�b[��j��(�i�dF�*��+��5S�I�	Y��	�����|�z���*T:�J��>�u�N��%z�Y�R�u��d �^�X��i:��CX<zӑ�%	I���{��E�ړ���C�]�rttD��e9�����<td3k�������j5䨣A��B�$I�9�P5]���wY�C��@��t��VJ�Y3TD�����0�4tߊ�^�6`/��4�w�=�����7㪀��8??���<<{opYk)�r����\���9Vf�~��̧��Uy4��vm]���Ȩt�A���~�7��Z�ӛ�9�S[�ڊ�j�:�X���n�g�"���,z1euӈ�׎�<6�ocW�-�I����+�CU�BԪ�B���j���X��Α
��bƝٔdS�%B�i`������f|�����͏Π�e�V�%V@�%;�3{��|��gte˪ڐs
R���.�v���k�z�?����7��}��z��?��˫i����)���t2�|�B%)]/[�Q�-I2b��#wB�A6�gPJ!<�c�h�r[qz��
M>�1���ts�k�z����ZۋPj޷r	X�K����]Կ���s��c�nv�	]���8��q8EPH!~���[6�m���c|.!D�g>Z<�bmMG!2_��?�eY3�r�1�����%e���l7�x�X	�Ƒ�m��ߴ�o*��c3�h��}���� ����^�3�4A%)�4�65]�q���n�v�Y>eW7�uM",Z*��"p-3�Х���,�ȲP��4�3�3zԃb�6�"�i(��=g)%H)Y]^���g�
�I����⌬mcd��Y��/�b�{O�S=z�v�9��2f��M8�y�����B�P��͈m+c~5z�!_~ݣ�i#�`|�譏�l�A���W � @!yT���׎�5��g���8�Ҷ�ڜv��,�ks�cLK^O篝��߮��l���,�hOS�O��G�ϱ�q{��Hb|}_��;ʃ8�1������q��8���UD돯?>Ɔ�e��ؖW4M�u32��Ɣ�ؚ�����R	Z��I����c��	w��6��K)���r��vO��}F��۔�X.��}dS*H�	��v�K�鄗/_�~��I�S��b>a��qw~��?���t��O?�W��3ں�b��'O��c�<D��:ö*YoK����sre�Z��-?��RJ��D���.>�A��]I����qw�s�����nKf,�S4��Bd���8GT�7����FD?j����1Pqq
�{�¿9yߠ�o
W�}o��[�x�A����5��c�4��{�ޓ �,碮�����$�f�mO�2z^����2v��H��G�{�w'�}���9n���p��=z|ȯ�~��b<޲%��I����y� QW�u��X,x}qΦ44�%�y�Y�� �y�}�v���y��{��̧�� pΑ�I���,�R��=�л^yF�7�LJ)doLD�޶m�L&ܹs�5_|�ŠP�e�l6���fP��<��~:3�c�P����WQ���cx�4�*�`�{�p{>)����>TH����rI�e���s.//)�|����iL����c�>�߱�=�$Q�؏SPt)���h
9�}U�1f�fn�ι�0����G%�Tk�PS?>�@ڵ�����·��7��so-�i�?���G�����6M��א��rfZ, �B��$H��iA����b5��!�׶����4��É�̪�搢���J���ל��p����'�n��))9=���Ǒ�i�q���=��]���NJ�	I:������BpD%�B�d��j��T�""�ho�l���O��~��S�Z?�& "�'b�~��=�Wt"����r��o����?������b�:�:%ܛ͆�o߱3������l�⫯������麞�X�QB�:�~�`]H��P��ǂ�?	��x�N85���H`�BI�s��=��ԑk��g��
qyA��E�)g�ϟ�� R���\8~�����^9���>MFH�I��sU���rz�؂�O��3v�xz����.��IEo��E�?�BI}DI{�A
T8?<��'ս�w�����.��3�8��N�š��� �v��r���y��7���'�z��@-��Cn>���]'i��������$Q$��0(��?m�N]�����r��ЬV+�<������;���i��������Ls���9;;�,�V�/����}��ݎ�,g��,˒vz�Zh���|���O�B O�d��X��D���2�-�!���D���e
�;li�9??g�^S�<^�l6s����2���&O��4Z��)`N#�� v�۶�g��9��x�IϠ:u܏�c��>8V������'���쉥��j'�5�o��#����~N�}z~O�����CJ�Ji��G)���DfJT�E�����ӱ����#�%!s����% P"K�*>�Nʴ?��	\���1�!ɔ��يZD����;�$���\a?�����a�s���:��6S$a��ǊU-	�W���|C\��O.ɫ��=P�9w��jA�l>\s�����Wx�怖��"]70���ȳ�Ff�s�x���al�O�ǎ�<���Y�!�$�C�3��*(�<#\��m�ɭ�OE��5�����>�G���.�SpΧ'�43��Fi�Og9/�i.~�}��ӯ������IH���O�2� -ND����N���i�t�J��1��lN@�'mT��rj_��|l�J��e�<I��L�A���Xq9�ϟ�K��������FG=���mo(�b���˳'�C����CL��JeB�c(�rnU+m��ir:+>^?ɸ���
!UU�Զ�������f3���*h
���v�9E�O��aX��<{��?���<ۗRryy�֚�m��,�����t�y۽
k|eYf�S�����xf߀�(8;;�C�4I�vt���|6.)˒��+B�}�v?�u��xF��$L�z�	O��{�p8$)�,c�\Ο����du���S��t��e9�pֱ�=���=��������fc�u$:�1�;��c����ܻ<Ð��)��D;~L������&r�5w�z������̿}�Gw�1����9�<<���	�W��R��i�"Q*��X���k�z;vf�Q��D 
��<�Y��mǰ� �C��6(�i����}0��}.�>�����-�O�H5��2X�S\=����{�v@>��I��\�k�O>w���M�_�P�P�����"/�!&��O��}s 
1V��Z����Zqڵ9Ţc��Ѵ-F)ʼ��r�������B@T��q�Ŀ�E����0�B�/<�ҟ�D�(�.y��7� SM�D����0�͈_@��G���AH5��Y\؍��N�c��kQ�̇� �C����jVIt����= u�ҋ�MA�t�!2�Y������m���ْ�v��H9rpǌ#�OZ�5ӗ�C*1���sŒ��O��B����w�)���p<yR�8
\D'p�E�/#�������>82k񡠍e�H��Z����R4&'�U�0;V*6�w�pݐ��Mv���B�>�� <�M���b��2��s����|�xA�7�ts�dF�VB�+T��n���
1
����Ȃ`]L����g<{��~x�ᚦiX�5�h���D�c��}ǳ/^�5o߾E�����%|�Lɮ��I�ZK�=�Cݦ�r�N�☌X���)���P�k�ՒLk��#���|ɛ��|��!-�"+	.���︾�]i�Jg� �ЃLꖹ��p�d-�����_���9ϟ?G*��(]˻����|D�t��,%��"[��*&F!R�&XO��d��-��[w!�u2�Ȥ��{��g,�˲���3�6�}��f���k�s��ۤO��4�Q#�"����2��~�)8��mRd�(�(P���§����������v�n�c3bL\H]m�s��8��֦5P&�D�@ʱ�vH�[m$���Ƨ���-en8;;�m[v��ܽ�B���j���~�΍˄��%"Q���8���"d$Sc4��x��~|��-Y��`��`ً	��D� �`�Xp��>M���N���d��j���t0��>���������_�������nC����k���^����P���ʒ����D	~��=e!qR���ap���;;
$�
t�ت]�}.Ǝ �o��x�D&�*PAPfi,�<�(�>u���H�y�n�˧
��t�:�Q@���X�%B�q��'n��+b�H�p� =�O+����)�\���S��Կ�T�Զ���㛥�+�?D9��� S�<΃���q��O��s���O/:fD�0���ܛE�V��ߝ���+�=l=O��p^��o�[�kECڐa�[���8�K��[����I�%��G�\��-�������  7FiD��3�$���B����d:#��*���Y����E�gS�����7��6x��TFq�S��\TX�ڢ��$y�R}����|���x�C����?p8�,�
��*��s���l�bU��������Ȋ��(fd5��W��
���������*LQ^s���H�T���V�(J���2/(2�s�7#��1�O.��mn�mE1V�	ў,E�X��u{"����.��n�Q@�ԋ����⼣\ԔՂ]������ ��a+\]=Ee%�M�,J��}@���ZCH=�ΈD���F#$)��HI|�!r�ӫ��ENf��s�CGP����Ue�}���O�KY�c����Z2�aE���N�j�ҽ��#f�L^�"~��֜]�s����_~Ż7o9�Ͽ��?~�>|@II>2(��y���B%Q=� �N���R+5�%H�˳5����ȹ8;�*�ѧa�1��_���")�B��(�L��H���Ǝmx�D	�Y�����u����	~@�i��"�[O�>��$�*�ϵ���܂�cҦ�$pgQd�E���G���Z̬DgHm��;Umw`�Y� �>&���Iϧj���v�2��CO�E82Z&|��7
%eB�>0�r���Ӹ!�ɜ�����(�]�����0�P�-Sw�4.?�0:����c��^��[�1��\nQ�Vq�Q���g�T�z�s)���z��"�}���N�瞟�J��oy_���Dfb)���U=�����=���{�~����
�z���URE���V�/���3�^� �'_�(]P�%w�->���n�<��O�;��x!0J�E}�>3e��E�9Y���)�B��Լ�<�������-��#O�gp|����Z$��I�|��е�Li
c�#=�ﱶ#��;g�%_����;����s�EN�$�9��#y�Q��[��з�0F�� �4]��5�1�RR�ת�9�-����R%��;Ye���������?"���n���X�ov��|Hݧ Z�0
��e��zEQ�l,1b�8���RbU��X�Q�%���<��ޠ���+$����Î��߲\�d�5��1Z�(xb��i�+�Qo[�#�_(9�� �$�)�A�D�ʪ�þ'S�e��v˷�~˾9��7ߠ�} �d�#���k�X�����1x7�W%"J��'Ø�Č0BS��%�w����3^VW�Z�.U��\��k��<�������j�G����Q2� R�A����X��<�zB���i�V�WWW����{g��"79�w��Î�*zB�۱�	nD��Hԉso��2������A�� V�{��c���n����1E�I��wAҁoۖ�^��9Ǣ�0#Pu�����A�H�z�=��P�����'vO ���[ i��u}L�8�N�&"͍�'����@��J�u6w�87��(���,�,��X2��$��	#%B&n��ux�R$�^Ge<<^���ؖ.�4/�G�" ��a�� ��d��g^<i>���M���3����tf��o��q���:·� ����8���cro�ı������{�8F"�Tm��,)��u�U�ruAY��E@U��9��!D��rB\��$ӆ��3���wI�.�ԺtCZ8���cۮ4�n��6Q'ѝuQ����o(T����|���l\J���x��!�Ty���/Q���x��g��-�fCUi��1��PXk�<���
޾~C����T������ժ��n����kt^!��h��<��b��$a�麎��6�I�Bf�\�##���lt�27,W%O��s��)���|�曯�b�7�v�m;v���kr�@�z�����v��nK;�/�<��ɓTኔ�<�<C�n�|؋"��E���g��5m߰��I�    IDAT�����"����]_�t��з�ဪ\�#W$âv�2b@��G�!xB𩲕*%��2�0 ��(��>�Ň��Z����?���i���-FJ��� ;@Ŀ#�'�<����".M �<7�9�%�ԉH���19W Q(#a eF���n7�=}�n�u�*K�5"˲J�S?P�@��;Bp�{����G��Z� ��� �,߬��oZ��-��~�d���n��m93XS�zg"�����0%�$4��Y��L��n@*IY֔�s�I�*A�%:�ġ'2Ȉ��FS�X���5�sk�õ�a���T��Z��=���o�b�Iv�(IQ%
�)��,+�q����jƮ�l2�
�0&Æ�@��Gz�z���2��Z�M���5�<i��`�$i�:�ps˅�uЊ�6�(�! pb~4�)p�;�����[�'�RL�lSz0�8�uR�z�ql�ρm���)(M�����z��'> 9����4��>6�wN3���?�R��Q�����+�O*������|E����kF���O,BL��Pd���j������/��/߲m�ed��jw��4�OT0)"��$�
.�I�97"K�=�㈴�3���������j������ih��������b����O(V޽yG����ޡ�d��yzy��YX���Ԋ�j��26�_|�����Bt��۷o8����;�0��"+T�'���+l����8g�H��m��̫�
�znnn�1Τs^UUzm�勗_��_S�m�#��~�r�p�YX�H���@�-gϞ���T�)%ϟ?e�^�;���{2-9[-X�u���[�11��z�.5�'�J7t��E�Q�o(�v���2��-W��|���?��SJv���.%y
��vO��M��T��(�)$�;��Ebj�y�����/xry��W����&U�.�td���W/������#.x2��YǄ�ȵA	������tm��ȄH�S�sBHP2����'���7-*
��[��xo����_%�����s��se���Q��`�/�Q�����a��4�_y�㇁�d��5/�>��rv�-�.�L��ȍ�|��סd����HqTn�F��6N��.M�W��0e��kYM㌁A��#� ���R|��yZ(���s]ؿ�3�ׇ�2�C<�ӭ�~�sꢌk�#�Y�7�v����wdy�$���Be�3cib�L�}3*K�fѤ8ƩS��I�I�#fz|g�3�)(�"��c܈�
�Bc��NZ�	�e<�(�8Ƙ��YV+���3�1��m��럔�� iG���1�	�k:���I}�����X�>�Z��Q
��^(����a���Av:I�]��'$�Hm�f/bő��R�?IV��}8�ꐜ~��{�������Kp-j����H3#7�3SP��=ϖ+�����[l�,//��P׆X�x�8��o����e�(;z��Gn{��p O//x���;v��g�y�R)����=����%������|���N2�Y��d���Cjwe�Y�'%e]�4�e��nOp���xv�@7���+����;�ίpC���ʄv�򫯸|�"��ƛ����,�ā�h�1R"F�	�wqqA���;���o_�4˲�IY���6?���|O�\s�Af��K7�z����3����n�qK�w3-Oˤ=`���b�1�E=K	!X����d{�'��/�'�!^����f�q�#��|$*�bU�����ï���w�azq΁M�kY&���H�������:���;����jVB��Wk�����k�4*,pqq����y��W繺�$�i뎦.��i��޿e�l��(�
�>
ھ�Ϣ�)��6�E]���s�a�w��{�CG��9Ϣ���7�P������,�
��d!��m�F#��YiY����B$fJ�kv�6xV˒�o�+2���ež>0����Z���?Φ8��TKp}�p�*Ό��Agj�
��:r�y��	O�>I�~��ȝe���D�V$ oL>�����Ed�<�����O[b�$=��L�vhx��-n���X�,��6�Q�J)���%?-�$
I���H阺����Ԏ�v��J�1<����FY�<���0mi�O�E��`ι�z��f3��i�t�S�ѡtԊ��ia�tk!g�)F��n����ݯ$9y���%ʓ��H;��J*�h��v��~I7zJ���x���X`�S����~����q 1ƣ�z(yXL�idq���'A�s�{��|��}�w����Bd<�#���73��[?`�E��p�~`0P�_B�Lv�mG׶�� 7�$Z��L��L2�������ݛ������ω��_�@�yυ
8;`t�e�)�{����&������j�eM�\pyy�:D�]C�Xt�Q�5e]%�5�ڶ�r͡�����.�`��c��������R�
�{��X�+��-W�s}�a�^S/�Lݯ</��Ͼe��RU9��z��EQ�㝯O�HE����6��#�7?Q�^���7x2a�MNq~���Sz�J���_����{=i$<C]�X�=�n'+�m�p�Xs�ZST%�U��yˇw���^�\��6A�Ed����%��+��>�n�*�ɓg<���_~�:8����ٷ�u�^�)�rxϻ#��HYs��j�ex���w��޼��H���.����_���Eśwo����<1t�sc���ٳ�o��z�$͡'FA?���$׊JI���^������QV�Ҵ{P�����_s��)?��EQ�o~�b����4͑G-R�?I�GӤ��z���N���p��*~��߲�n���G6��g���%Jg\>�BJ���7�gg<{�$����]�ь��j�b�\�FMӬxU���+���ӧ\\��ز����z�Fk&���I�7�|���T�=�r�u�_��O��QR��Fѣ�d�>o�\�v�0i���z�&:�P�;%��US�ͺ#�&�>3졪��z�����u0�<���~�<
fCZ��e?���J�&��j���b����<�[OZ����OO':;B���d&Қ�?or�+��n����k!=�����^P�2�������X,�jֻ���R�cc��Iʣ3�������ɩz����G�:6Y)�Y���L�{z�'W��8�i7��st�\2���XNя�$km�
��bbH��1���q~~�y�$6-?����޼�28�`�C��z�y�B�KI�3�b�`A��sr}}���ٚfբ��:����@���E�T5��c������޿���/�5[1к��2�U�*�j��EQ��%���r����^���O�<��ũ6�1�K��`ɂ��yǫo������*D���%EV|dQ/8;?����o�������ʲDZx��a08�ɲ|v�+�+L�t��������O�?|�%0���9�,��d�S��Q�����/.@H^�z�0)iv��D��0x8�\�H�0eF@q��⃥4
�5o^��=��{�p,��8	�,0��&7�i�ϟP�lO����#�K���h�~Ƅ,�+B�#�9GɌap�Fh�"���w~����{����xvqΝ���bU��_Jq��)�V�=-�E;+���B��K�H�=�f���O����~{�`;2�����_����������~��@*�)rno�o z�?ί�k�|�x�I�@k���;�L���咾��$OJ��I~9%$z\�_��W�ݿ������{���r)~������&�G�@!Fa�������l����]�G��8� LB�Ǐ����@����B��<�!��1G��S��)��c ��}SAx�2�W�D�̔���Oz!$����1j��d��t=�h��y�Zb�Z��.nR�9n� �f0޴io2���@�����1��] ��y�>�n"9ʿ�(r!���=�d��@H}O���7Y�=��ߓ���4��w^@g�	�B�T��(�BM�c0Si��l$��w;�PR����n^G�H)t�}� |!�i�y�ƘQp�xbF�I�>E��.�OզG%�1$Џ�C�08jY���#��CE���s~���/\��=�~x:�~K�O��u7˺J���a�'x�B B$���LK$����n���l�4" c�}�\�# ��nߧ����țw�X�V:�����'Ijr���h�0@�(c�U�:�v{��f�p������D�8�:7�h��w�Wĥ��f��h�pm��M�P�e��#�/�>��緔�ݡ��%���\���w��l凞���]T#�1C�Y^�B�����	�7\��Ø42����0J MF4���G��eF�٧žu��F�=û-ݫWd��Ry��MVB�)��˺`U�4���~�P��b���}� D$x�r�B/+�N�.�I���Ŕ���IMyVSE����c�������.����T�fY,h������%��բ��r��z��Ő�v�&��#Y��H������e�Ѡ�C�;��翧{���]�k�+�}Ca���_�Ǜ-NJ�q��	eY��Ke�ú�_�G�I�iD��~ٶ=]�PJcjC�"��5K�����?������`��g\>Y��w�,oO����K�4%�v\^^"Cd�%N�p-eA_*��Fd���]�&�H��z�����-f�q���z�տ���O����f˹
mK��y���.�EDͤ�	�&c�	��4Dy�C0�_�]�8��u�m
BTD
\�z��F���]
�X5���H�s�vkq����$Z�f�|��J��J�R5*��O
z
���	Kd`8@�c�/P2'�%�.l�B*��8���P�(}�tY�aSI�iB�G'�!
�PG	\9�Tg��� =��F�G��8���������L������L��ᨵ=��O]H����c	59��S�ϩ��)�����?�M��Y�rB�q|�T��<Ip�/I�	�4�9���o)A8Fĳ<B�D9�\��2��|��7<��oEI�Vt!��n�l3ue�>e�Z���b$�#�	@i���(!��}�[T�(�~ ����*Bi腤�
'E""���a=&+'ZgĶ�	�.�U��O���~�Ѓ0+�s�
%Z+�"��M������r���cK0F?zzK�.���ؠ6}�m52BH�!8Ę0˳����w,��L��.OV�=�W�m���5r�γ���U�r�@E�W��48��n6����'gxgi6w�-n�qEN^�dv,E�	*c��s�Z^����O��ف2�i����Mߡ�$�9��	�t�88ǻ�{}���!e4·$��<C�z�^*J�!n>p��`�z����ۄ�X�hchE��9����{�X�q��v�bn?�[�=����}���������l��ʜJ�b��D?ܱyw T���*�ȃ�>PfyZ�"/R�NW�uD�~��R�+	�;�?~�v���Z��P�M�A�v���x���{��s�4�egm*�LF��m۱�5�p�q��YGPՃ��̐Z�h�6|K��p��>�r�#���"�1H܀9�P�5.rR�?5>����/uh�����A�|FDj��
�:+(u���u�CQ�8g�CwoߥL3y8j�8g���ּ|�_}�BX޼~���5�����*tÀ̊�}YV�eYf�d��<�����R�d�!��F�n��x\�>��\-z�"nc�{�ܜT�S�KU:����� ���c��'�q��1 �����N_{�B�o�c�������E��epq��N���?��L�tOM+�����R�h���(�9X�V�
M�  �zfs<MI�C$��x&�U�NZ����(ȍ���9p�I�Vl)	y�I�.JE5x�j���(?L�=vi��QL�E!e�@
2����Q� 	����<����I���Gl�!�;�,Ǚ�dZ����D�8+M9?�?р���%}�f����M�/P"�o���Gf9�u�S�d	��ԩ#��d�	����>I��1:����>$��R�];�'�"����w� -F*D�ئ���?X`�/������=`�.%>���g+@��){nH��0 �L�4��k2TY����ha�xv��129������->�\c%Fns��H��M��)��kJ%p���-Jex�#��r�jEP��}��05qta;�mO^f��ι$�;XLYQ��X,dJ��;��+��Ƿ=��ےg+4���i�޾%�{��s��`��e��|C?�L�{!�I؈I��A���1�Dl�}JB��)�ŷ��jQ ���J"H��|}u�~�s��{~�����T���*	$�f״h��)M��0�N�:�8{<���t��@��O�(�5}�ɧ^���PH�,
�В�O���YE����SA��݄�(�pD��Y�����N��aF���x:L���K<Iv_^^���6��<}v�bYqssû��]�$�6�0&9�$|�"+���_�����-M�p��~������W*@����O����Dd��������#'Ú��>�{""���I�Q���F0���|����\?3���cB�Rg��8'ѱGj��}���R�s�AN��.�����n���T��w;&���4H$J�Ols���KJZ�}#ƈ�728S!�8�(��\h�����w���ӧ\>�;���[��
ʺBGE�m�a�$Jy3�qdڻ�>�T9/�]��7=Uf�lr��c�l�BV%:ϰB��DgѡG7� H�NҠ�Y& T�$�v�
ee���J�� )�Ż��ɤ8�H�Z���bH��A;�tj7g#Z��Ĥ�d:�;-8��C(9���vD:?	���*%��'�a?��]���a 1F!�D�>\
^1K�5�#qp�h|�(����ua�T���Nx�Dy^�l�IH*b�
;*�%ݟHt��e$�\�GhŪ^��O��b��n��-e�@�K���:I`�n��%#��q.)�V'�#C�.KL��G�2��{޾zGw��H�Pg��H�$�|���J%^�H�͝�lX�%a8�D���!�Hbp�C�Qf��k�����^R�lc�4�sm�x����q8�c|�5�<�w=28��a�#[_�:���#�:�?[����(ߣ��`[D�	>�i[ľI�����`B���21��wtCK��2X�@eJ��:������8�ܐp�|H�c<���2x�~>D>�>�p�\����}P�Lq��HP�h��@� �'�[�PdB�뾐z�)4Bl��s1��I]Zk-�޽#2���R�u��~��-}{���JM�7I��;��EA��,�4x��-�zn�����.�ĭ��T�ਥ��0��3��~}߈�Է$Iת �Z�zq�_9�'xz�sw��	�@M �����CO�4N?���x�&���gH�Н�L�J��&�od�D��L�^�B��	�%"���6�+�S�jq�>N؉�=��!�y)%(K�I�L(�!ۆ7�����p�����kZ��Y,�i�v���g��ClAILV���A��SK3+R���)F�,ݡ�kZ����)@ .&\E�,�Li�32V�I�_�8��W��>[�^�1H���[�߿N"0W/8��`}~�P������i/�i�BQ�Q3FT�	�"��}��s�0���:�6��o����7 �&���B��J9����Y���,G ����� ��F����J���D�@h�}�� e$��ɲ^�EƦ 慤��G�i)�2��]��ݎ	)�D���)0��2cYVܺ�E�5����GK��*�z�T�4Jg�F���p� ����-�0Q"���mQJ��Ib���*�*���kpْ�fOU\\=	���XԈޑi=+�y!`ԑ��"�ĈC ӆ�6H-\ a��=E���^�4�Pr����혋,�u -�*7�v`�6Ib蛖**�U(����@�8�������o�w�sM�5m��}��"��DQ%-ߵ���2�ʳx���46�QBY�4�[�0�g�    IDAT3�@�>��j��Q��\�9{vž.8�6h����p@e�4<�KS3ƹ������<�[=��?�p�
e�p�	�$����ij�O�,��B<��pGzm^Į��јhZ�E+����}��^^����-W\__'/�U=v�����|��w�����g�5�g���)\;*�XԆx�+!�b��E�؁�
�8��#�?i�ǹp\��b��Kv��n��G��G����
!<ʕ�S'yZ(?�����#�b4���Ǆ��q�>�D<N�O'`��?�-B$:Z�'�C�"|?��G����5�Y�d�c>��y9-qܤ8L$�If4Y�	~H��Y��������g0��}ö0Y�,���Ǻ.U6JF�JВ $�;T�}�:@�����K�^�Kp��Y���ĔrnA1��'s!"߮��e�\�*
��)E�q;�D%.�n+�m����J�ȩ57�"H�p�$&/�C�pq��Z�29RjI�
���W��$�9�s�������e�Q
;�H�Uթ:��e�2C��cBߚz���BI��a���F�e	|iV��Ւ��6Y���EU�I���l���x/�ă�<O8��Z�9f&�&\�
@����UM^e�,r�=���(*d =&J���d�|�I�%�5�v���uQ�X)�G%��d.���˹��`ڌ`#��Ҭ��(��܀�t�M+�z�(���O��3C�B�������=�YK)��
�Ck���u�4-��F-����UF�^R,jBL������A�����.�q�`�.-�q���/��V4�E
M.�vH#q10DO�T�R�ZKZ<K��L�M(�?r�s���,���>�mZ��k��=?���mG�e�<��8x*��Y��M�lZ{��sA���>��sa(}XIP�P
i2�R&�X�e���*#�KI��1��xR�K���9�6�<)�u]�܄�+6�-���,�ɹ�<�d���������^5`H����ݖ�O��XV����@&V���gf��a�|%&[1B�@8s�?p���A&���gH��5G1
�L��Qs�>��Lx|�s3��z>�h����cHf���Ǧ*�~�`�v�i���H�����9�iw��.�C����Eʔm�󑺗�<�4��� �܇���@JʴȐ��O���*c�]ϡ�� ��� �O3HQhd�,U4n����.D�c��H�[��cbt�RYf�|�D��EGoJ����@jOm��t���p׶i������FQ��Z
���-��~p�(�$
��9�G�)F1��|q@d�aT�#�a�@4?X�Ц�p1�p�p��d��O�	��E����|N�ԝ��m1%e!Ң�(�S�5T]aQ����U�,�*d�~�cp=}����0}O�#cю?� �#F'����,Q��B����dJ�L�ƬWp�DW�͆���A NXV�O��c�SIo��5&*$*]�UAY����xK��eIV�x!�%.�;�w{D����;˻��|U��UdT�����z���<�w]�,oP�$�A4"E��ZR��{:���LD�?�41�ѭhif$5�[�@R�%�� P�d���m�a�sMV�fbNDFf�{3�ۭ����o�ʊj��U�"㐧����UQU�ppZ^')E�����GYv��,s�D"\L��!�5�8��e��g<����H)�u[���.&�E'�l�P1�V,t3 h�[�2BF/�N�q�Pq�qa8�����"q�b4��ol`+�j�$�����GY\Z�r�ݻ�TyI�Ӣ�����{;��b���G��k�z���[.��Ǵ{	F
li����ե��:x/������7��`�����h��z;�����')��j�]�eY�����eq����6F��%�2��6y��j�H=��h�G�?�����٦���^X�����+�����W�=�"���	�����Z]��Q�j���%%�Mm��>E�QW#���٤�'	��~b���	<_�B5A-y�|��4����#���?i�h����A5k�3)�)�`Z�1K���_S�7�J�>�ɹ��W�L��{��V;t�'��LSeY��1��X��e� S?$xuA�n�n����q�������V�KUz��-�k�j�j�9���� RH-�D���\�*�ZF���2	�Fh	"x��:��Y��c
�x�0*���I���]�X���16���A�e�����S����j2���D�Di��o,�,��5�JXЮ�\�7��tD:����w��b]�_��"/,JJ`E O��`DIU�y�\�I��J��D"8t��YhSjm�nD�mK�0��f+���YCUYzB����ʃ�>������L�C��ݍ}nݾFK��W?��^a������%�#<�i��?�N�l�k�8"mQ�6�ģ��*�/�h�.s��md��~�U�т��"Vt�������p���78�7@Z��	2���@hG�%v�v�P��cd�2.=�јq9�{�T�SN�-�iI�~>�K7��+�-�P�*��1�8����ҁN"��I�WZ��-E^�������,�0��WM�X�n��R8oHZ��������ۣ�=�xD/k3��Jb�Q�$m�Q#V�$C��sZiF�2��Š̩\A�vY<�B����T�{$B���������5:+���o�S6jm�$!�(�H-��)*��2�I��,��9��u��I���>g������xʎ���f������"���o����a}�7%FJ��3���xmF�qT�ϛ���i���y�#��,U���K��q���2F��lo�2�X]_��ɓt{�9q���P9�B��5�L�����q��o���F�uV[���M��[<7�އ�2tKJ��J�w!)}��80�Bq�C�i�� �������P*�51������AY!��/QR�$����ak�HM� ��6�CsI�xc��T��)�.���8wo�*��̥D͂�I�����l�ڡ[�$'����msJ�P����z}�@���k��7� )FX��v��0VR1����QM��X*��9�iD$[G;�I{�E����2ma�%FÊ��1he�o�!�cRgIDF9tdQ��Fz��Px�phZƓh�� ��}XORJd�#�����bhF����ᇻ����Ŧ-q��EF�\Tx$RH��n���K�s[�07B�+O���e�L�T	��@DF���a��evF9ى%�#!�%#�B����bm!���g��%V��3V+D�%MR
�q�N ��)AA��#�@CoM�G★V���{����5��1z+,w��w�����e���ڙ3D������sEp��
kw�8�Ne��@)O�@��� I$x�x<���_�ȓ�Q��ʋ�G��"�E��t���{<�{���3�s��7����W:;�N��YF�.��DB�I,)���/�h_���a���2�E`�c*"_Q��X_]�n>������T&�	Z�����Gh�I����6��sh�;)��X�9��&�z�ÊV'���[2N�R�Q�-���8��X��v��xwD�#���}I�UUn�j?
��TD�B���CZh�\os���tD;Ѩ�3Ғr[!UF���v��mR4�wB�hLU�(�'�<�i�Z'cW�$���n�#�����'�S �����ї��5	�&�j�g~��ڭ�'s�����j��Z(*d�ֱ�ft�k�K�qL0��N��kȴ@*(�q(�E1�JQcFň7���رc<��3��x�A�w+��<����k��X)Y\\b��qt�����x0��<���pQ���"���Cð��bLEP������N>��
R/q�B)MQ:��T;C�b�ILUxr�k���g��I�6��2�wlY�p4=9J�f^�zpj<|��;��[�����<� <8�Q+�52l�,J�:���Q�{��T��V:�����L���ｌ1!�R
Q+�5d���h�9��G q�缴��gS!��k�����Ц�
�7%N"�w���b�����s<��o��+?����B��-����E�>�0�w^���RUȎ�Wo�{�$4��4��pΫ��F�V%�?���"��apa@�I�C��ae�5�ʃp�`Y�T�M"�T��($B
S��&]�̃$�"'��ưr�3<���9�'�K�6�����Ȩ�eū?����]�q5�۪ڋo��iw_wsI%%Z*��*K����|t�6��n��"�ݸ���E����}g8��Ctϝ��#�/=�߽�ۺ����o�H��(k�T8y��$*�q�e8��=����?v�ň��ȫ!������SDKQ�l�4Y�ȉ��$�k)�� ��4����"�C� ��eA^TT.(�	�ϻ�����"G��TN2�-�HA�(Jq�T��ri��GqPī9Z��6p�0�Ag����ʁ�,,D�H�Jb�O�ΓJ�U�Mק��I��N��-�H"�blU�i���^NH��D����r��(�q֒X����8Y�FY��
OE���ȥ��%Oe��ֶ" $�!�G�y1�ٳ� L�D������r5���'{���J)��Ⱥ��Wj� �����!�~�v;@�EQ *;-�% �y�c�r�u߈�^��`�ݻw�~�:'N�@JI����i�q�]����&�N���ʂra��x0dow�*/H����*G�!�2.\���k7h��t�ݩd��C�b7q�xF��I@	P�bX	�DMI�q�I��`#���������v�L!��Η��Mpc �B8h@���[��d����>��z�u
�;��1��s)���8R:��t���{7�ɯ!&�����Y;Z�~������qk��i� x^N������|5*����q���y����������a**c�(��������ѧ�yύ�����TÄmRB��?j�_�8���h�\^�F1&��:������$�T;�&�W!��Ř�$×U@�����.�@�Ҙ�Ԇz�L6
[�X#:K<��Wy�+/�vd������&c����j�&�ԣ�����������ڈ)!�5qH	ХF���fQB��"R`��,G�����|���]���u��i.���>�W���ĉs'h���sA���6xQ;�Anb)P��z� �뱅�,J����ezkk���9�����?�H5�8�9���(�
IYI�B��c�91�!eh7k} �� q]���}U��t�q
��xDG��`��2g1��k` ZDآ�G)cgȫ�$��YJgơjxS֬;a}��"$�n��j8��!�R�2$qF����9[��T
��15+������2�X�o��U��޷��+���BĬ�Cai��a�P�v����xD�Gc)��W)5�U($V�EI�b�uӱpJK�Wz�Lg�������7�?gϡ���~��� �9#u����S �ʗ�D7z�_��lS��3h�J+h�;�T��}PG�~8�I�$	����h�`0����:����]��鰼����uN;�~S+͸2lllp��e�ܹC��bqqqb��p"��օ����4q�a�������B'FS�����65����9��ƙ&<od������vMny~�挤�e�7?�k('0���{o����)��>x=�:��򽾑�UQ�u+S�����5{�}�?�B��ש����j&I1i�1�H4���g������߃�Tã�����9���t��C��w>Tg�������
������[�E	�p��#��|��k��u�=� <�,��-娏��z�C@R�M�?������D� ����Ho�A����3�nJc�Vڦo�@���������;Ո��Iu���oާrA�p|��asi�N�uđ���c���p�_�����_�7Q��_�q�����'��,��Os!�"�!�K!��Tq-)c1am'��J2ݡ�$�b�r��ϑ��Xai[�͛���L`h�F�ȲEO� �S��ȁF�^*��vn�@�n�b(�
)b�mk�/�-w�����1B+>H/�\E��_��9�zF�����$g-�*1J�@8I�[ʲ
��D-T����Dʜ����9Iyw�b�@�N��UCk�u9nu������77�mz��i�&P��S^���g��d1�x�#G(R�mc�C���,i�:�V`"���ʖ,ʘ�;D5�iJ�t�瘟:�2�hyDh`��9RT����$!w��bLi�TU�CuJ�j�!:V8�J��P���@�yo͓�8��\�Zin��YsJ�Clƿ4�?,=�I)������	�o�D3%�ӡM����(�pv>���N������G�j���v%������.ֆs��V��Ͷ(���a������i�P�<��>�n�
x��nO�i��+u��=9x)���u���[xaR���M��m��:��u��	d�|�ɑ49� 1P�>-�����C�����������+PZ�肝ԛ�P�@3"��O)%�����><&�r���:g�'?�O]�F�9P��'e���r!���QS�јx�30�!c9{��0�[ ��f�z�m�ֻ�r�i4��t�a��)����ѯ���҇�ƒ}
�W[�F���oxkT�[�ɖzTJɔ�����q;�Z�>̃G�R5v?MJ$t[�1�4��"�{�q����>��VFH��UYҎ4��.��������k�"I�	��Q��>�%����j�uF�@�Z2p#N["Yi��q��~�c������Bۈ��/s���x��G(��
0xT�� غ�;�e<�&M�'=@�L�!�lm�p������-sَ��9q1������-�FG��>1�q�;�u�b-�"�N$�P�o\P���
����{l쎸��{��?`��-.����]"��Q�"%ZY���'<��/r���q�V�%,�ek��5N*Jk� �,Q2��\US���Bp���?�s�ݼÛ���d5,A�n !;w����8z�(~�>��U�qe@jA/!�N�q��CJ�Z�D�XI��\%ة`����N���S���y>|��<�ه��=�¸,l�w�2��-��5��;9ǌn3]w��$A0)� D�q�����)B%��~�yBE
k�Yb��J�-r�m�p�����g�l�zc�E�jU���>�g͡�����>����(��}8j�SX�:�Z!�ʔ�vV��i-۴ߝ=��(BɈNw��]�@�N�h4�/r��-��sb��jF���$�zR���c�]���۷C �LhJh�n�iy�#����(�����^*b�pDQT�Ee�-.��Qpb�)o,��K���qu>1e�`�N܈���v�������و~Ɠ<tB-���O���$��Ɠ��C+�|��R�R�0�ќ N��aq�w�>>���@K3�`6�(%5��VL6��s������}~vτ���s������ԂC��Pf`�z��Di���n�.�Q�=ZH��w�wvI�U�������ܸ�jKF����ٴu��j�	�St��gL��u�b(}`����V�@j�^<��~C/[`7Ӭ�����LU��)��ݼB�y��Z����I}�T�fc�dQj B	d��qA"5/���]��G�@e�s�r,��DUF�������1hE��D�1g-�Me�E�vj�R$Bȩ�pd�ܘW.a�,q���ֱU�!��TJ�8#Z^a��yq��͋�e��^C�GJ�*h,(�fU݃a0֪}��q�"6�i���7���O��YK3��R���m7f$*���2��![ﾅ�Pnl�����C��Aǻ,m]c| -Vc\��9O�_���>�ay?ɱW.�H�0��x���SϾ���K���:_�+���u�R�ڙ�{]��"��밭L�����I�s_�=���;>~�"�Ns��ɣ�=�ʑe�������_��+?5l^������4mE��Ht�ypU�{u��Z`��J+&Y\a�"�E�PjTo���fw�#jEZ    IDAT�V�8�$�M>ܣ��Բ5iLU��\$8�WKQ�4q{>�rΓ ����１��ʹtf���r&Ⱥ������؄K0�xCEI�iVG�9S���D�SUU7gT/�Q�,��8�����7n�@�P�_�%� 7@ȿ�x�K��"�Cka8�&$��dúo��6R�͙������j�{�R�TGEE9������ڲY�\�)� �� ��L}��NZM`�zJ���M�$ 發�a��?��_e�� ����:@���}*t��Ej|�5^�a������î�=>6{��fU��o����g������BqP����|�λ���=�-q��	��V���Ўӵ3������G$+��z]��;�P:�������K�B)�	hI^yJk*Ԟ�=B�%j���t��*���o~̛��;�}��v�ۦ��qB�<�Q�����,E��2�1�8�56`]ȿ���]��Ό��b�,i%1�0d.b_���kl,� U��PF�X9���H����H��0�<�|U��P+dDef�}N棾/'=��s��Wpm�g�~����#��n�~�+�
p7�p嵷�z�cZ|(GHI$%J� Z�@H�sWƅ!�8�FA\ԃ�T������X�u�߽Kn*�KO���,�bd���*��ǗYW�Vѩ����:��P�,Un��4�lt&�����l|�>�����?�3�~��,$�����ҥz�>���<���]��/��{�9�.K�8Վ��:!�` A�JȺy�����u���u��XLڼ���{x�_�ܳO!���_?O�����Ӝ}�i�`�wo���1���\������	�%�DctD��gx����!f0&����죅��Go���w�Ӯ�~�Y���R���܇dT��ٓn��y�~�!l��]���P�!����-��Ҩ:b��j�'t���U]m>��[r[��`�~4�؊$�a���,.��j�fZ�Navc���T]�i�Y]Me��-.��N���;&-�a0p���~*��I�%���zU��b��'�w`�$�VUh�2�N�I�%���,T3U��`���f!������S� ����r5iB�eq�Ry�Dk^(EN8;��w0��׀޻�g��f�f_�@��y�4j�N�|�>�\xp���N{�/?i���~oJe|S!����j�yB(�^��ps���O>�<��p���b\�:���q�|�%�SG�_~�ŴM!v�bX�v+!V!�T:���`���҇�mv�M~�|�)= �#��7/q��Y�d~�}�Ɣ��!���(�G$$A"G��c�*��k�{�2�t�İCZ�E����wٿ���[|�k���ˬل�)�*�|�e�%-�Ȳ $Y��׈��UB��f�R�'N@�S��l|�.o�nr��N�y��J�E��x���y����,u���o��bx!C��H� N8���r��� ��f5�����.wy�gy��_A����k�����o�	'�}�������[����F��e����Kʪ�)��T����i�mr7�g�O(C�;�EM)J.��c�S�������|�����3��x�k����|�k��x;��{R#A��9Lc|�|MUպ�cL�E�hU���.������8��s�G��%$��!KRį��{,?œ�m�{�G�E��3�D���g,KKt�1
lu�|�¹G���v[ܢ���R|�����e�jĊ���z�mZ2"���5�0�`gγ�;��8��<��O�>)��}~�{3���� �:�����zj"#���s3��~"��@�B�:/����u�]�B?���WB��������q��n�)˒��� ��5l�	scs3H�ַ��?]C�Sv}X�q�T�b��o�ck��8A��xBC�	�M�� �|~�4Z�8Ϟ�$B���c}�����ZX�z7!��=^�Щ5g@C�l�l5	���.�U+��p����`N>��SI�ۦ��Cɰ?` E�+���`��-�>�y_�wCl9��&9�z���4BW��F�>j �iޥ!����MbŽ9l�tS6Z��;,��R��� ��Xh�����!��DMJ�П�	pO'Q\>�6���>���=����N��vA�CE�*=q�M�nS���n�l�lӖ��(R-���=�8��ȇ9���شc�"�����@H��aQ���qn����o`���+�ݒ�^�m�EKf��m�q�4P{yA�3d-Ϭt�D`�z<�����`Y���.�l�X�ٺ�7��O~�9v�$�.Y,aP�D��CW�d�����%D�N�����Z��c<��B�0,�(����y�%IG�G����z�W���=bi�a,�Of,/���"�Wo0z����"V�ω#E"%��(�TJ2J���
mJI9�Qv.<QǓ$r�,��ѿ%ZiQ?��3d/<�����C��n��Ǿ�Mn��Gl�����)4��P�*l)�S
�5�8�����q�BR(O�-x��gп��_�K��N�%:z�߾�}��`���K��q�]���DI��P�D��	�g�vE�$�D�@�	��pP1�\�ӌ7�)�6ؿ}��Sg����*��#]67.����� ��.E$�s�V0�3G�-�ǎ�$Q��	IK!}NY���|���+�}�[wn��?~��k�1�����I֏��+'��'��9���0����"'�Q�
_��%�P���ǁ���CK�@�(%�&�W!%B5�k;	$!�?��Y���&ha�L�5o���.�}�(�/عu�U�`� �F����)t�����q[d���U�j�xc1U��Y�h��J�,΁��(-Y\\dЧ��`��bT�y.��V�HMȽ���Hy�-J���(BJE%�=����ߣ�͐��A� dFYT���۪D��-�@����#b��R�L9b�����TE�":x�_�7���a����&�3!�zj~*��9:�s��X{o�:�����;lll��^dJLɁ:���k&0�����{�@���ڃ�~�L�3���=��j6���(�a=�?	I��O�,A�m�7$���N%��q�4��l���_�ƫ��sf��^��lc��������l�s�|�!��|�? �̼��<�?,I�b=�	����fh޻�������B��m����k�ȅ��צ_�ĺ͎W��%�G������,+�{X�2&铙T���$��q��{�nEU�Q�0ܮx�g����=ZkK�:)%1^	����cW@���O����T$Z�Т6�����Z��i���%���±��gx�+��������E�t�'^�gϜFZO����?��������H��Am˺����3��)5N��d�
�!"n����2��;��׌v�y�[��-q��Uv/_��V�;�#>B�q�߼�.�"����e�p�Or�Ɣ�s����ƣh��}D�M|l�;���m��K�je<�䣼u�=�����G�z
ٍ��;$�@G���QxbRG$Q:ja�8���Z`e�)M�*rC����g��O�u�Dm�5#Vz-�ύ�-�k���q�E�C�38������뤴dƸ3.r��B��Jz|��.����?����=�E^r�4}�E�Y��=F���J*gC�d^g)�21k��'�#4�m�ZjP����f��)��E:'�"DE�����N�[?�>f��j[72�UB���:���@x�T�p��9�iPf�:�֚(������ ��Z!o�ki;K)�b��([s�Ҵ�qMT��Ji������*Y[[����p��vw�'�cʰV�r@c�Vb��(�1�ڛ������\���U�'v0'욨�~���:��'M�'M�$�?#�כ�'��5����.Uk��	��l��|`=7�Ygc�}l�*���o�����c3�:�ws<���P� ��*�C��S ~�5^O����C�������_=���}OwZ\�v�wG9�}M��Ak�"֊Q���^f�V�V��������%����=�I���dۖH/�X��4	���%���
�'á$<8���$��|�A���3�W�q��B��K��Ω�����ӨXq�W���kT�1�Qv���}]_��٨aV�p�В�n�QY���6�ޥ���L��,PY�%�
K\�cܝ�@
B4u\ �?�ta��_p�B١s �"���{���?�"����6����ǋ��׬��8g��QV�e+r;f����������� �Y��b�n�h*�n�,EP��DL���5�����q��(q��I���;���嗹��5���,?�7�F���������� ��A��A�}���	�	�D�pV�ȓ���7��Xj�Г��d+�,9�W��䗟C�<EY���~����Ur2�Z��ڠ�G* ���Պ�ð,)
��i)ؽ{�+�>ʹ��S�Z0���o�a1j���ϰv�8�t�o�A�mM���56�rJ�TQ*�j�p��_x�Y�v�2:R�*$q�d)�;��9�ŏ>�oG��!G,q��p�S�N�Ѐ�M���z�������P��a���YƁ���-�_����6��������A�	�|z #�D��4���׺��ژ7n�sQUeY��������EFGh)W�j�|c�[i���F?R�$I%Rjt�T�5Q9O9
mj�3H��$	�n]���� ��3ܓ}Z�*������^���p�&����I��j8�S'W���i �������_��O#��^��A�Om��RAך�hZJt�911�A�|�>L�r��dj�m�13�����3�4M��%�P����']�����pXl2�p
����
b�����;����}=^������YF��%[wn�}�4O���uw����5��>-ie	EaqR�d��Z��'����(��V��O�q���H�U��Ǟ��/}���?�M�����y���d��3�G���������`4��A��Ha��q�]�>x��!R=be���x�˿ϓ�G���{�%	��*��;�ΠZ
F#�������h�OUUd*BjT����`�B��@ �㜸��������eƕ7�g�=��S����?ύ��om��:�˜���l]�����3���{�qEY�����a���"(�#[貾�N��E�t�/�G��p��!Y��������H����Z1,��y������� .����Fdd�=� �{���KM�Z;��H�O,�:q?.2�����?����|TW���s��@B�J�"+Z�Z%�3(KF��z�R��������_��ٗ~�����+�IU�͟��k�z���x�K��/������x���>:	��򯟞-RJ���z�"EᡨRZRgQ#C���Y�qe�:�)0:��.��_�3o_�Ɖ��?�*�v�ؔt��!v�::|�0�u�U���a���~�힛�YGA��}hϞ?��3*<�����~����_!�Q��a����_Q9�h�`4��9�1�n'a��CUU$I����K��I0��S2_�$$Q�I����uEK��"���!���Gv}�����w�ܭ�%�·�R=Z*��H��&�~��Df��%�	!��Դ:�ׂ�!t�M�{)T?�r�L��榓.g��~��E�3��y��u��1A�Jb�Z�l��V*�W����D����+W�[�Y��>��)���&F�NY\�=�Þ�����Ĭ1f:n|�b����s�8[�{��ɓ1���4��[�=���K<��SE#~�ӟ0v� �V[��i��W�.GD�En���wwH��(+��tT���[�%�z�����J9���fE��c�(�\�׎����,�� �C��'JZ<��K�}�I;X*v7�8�~��/}�;|���;���n �/�s�mMnd:�I0��Q�q�ދ�ng��~�\�@7����UN������a�
[�/5�)�7�S73^������%N>�e����.���� ���/}�B���?�g�,,.���kN_��+������Vƹ!H��p0w0�Gx!b���`gYZ����:k���E�-�h�ͭ�,�;G�����1���x�$Bi��':�Ig���s�*�T�巯��0NXH,$B069��%l^���de�����x��^A�MBs"B�DI�Xz/y��|�yQ2�,�p�	!p�U���k�����͎p��9�,����{�ט�;���^����)�kwXZ^
�3�:+ڤ��x�)"�X)(��b�7��O^f��$���=���}Ȳ��]����,�X��������cL:�ٲoqZ�I᪡|_�|���)���MX����ΩY���ο�j��Hش���bA%��B� �sO��^/ �P::�Y���u��D}F<�׎_�g��	`-q4e��1ιI��$I8z�(=� �~�������
�*�Cloow���^Y��H��L$i�ی��	c?M[��^Δ!xl�Fe��j4�.�fޞ4��dCMG}�PS�٣�7��䋉1������I�;�gZO�a��r�Io��(6�)x!'�҈܄��N��B���f)X�ZJ�L��a�L�V����n��O��nλm��It/�}<h�����|�0γ�^�`�9�j�)�9������73��)DM�s�}�D<�#O>͓��X8r�ko�����He�$������k��=��jBl�?�9��-"!P���r���GF6�u�X�8C���q��y�c.�����N.�̃��_����s����<��o�����R�+Bn���'*\�d�s(��{�]'����]��������dLe!���.�>�/|�ENY��y�������K�!��oeU"���)>D�k0�FH*A)$��%Z�#��=��2V�d�侵6��|�1���7����"E��
��x'(�9�Q^|M^d,�� �37k�9A�b��❟���'Y;}��^���Čr�tȻ�>"Z_�?�W,=�z�i�����D�U��;�>���tO��Y8u�~��c����w�����,�8AT���@K�rN8�:�,�Qc�ƻ,�X����ꔠ�!��(�[8gQq���Wyaq"(
!�ƒ���$&V��m6�����'YV����Hv���-���%n�_�;�_�)G<��9�.����~�)�1<Y,��1��a�3�ttF�s����/摧��K��C?.��DG1>��?y���m�o�`1ˈ���	M�5���:O��a�'2�t͞�R�,j�ݔ����v�b;�"�,+t+��{�hҞ!X�Eq�F�����Z�J"@����]�u ��%yYM�eA6��U��v��YXZa��F�����n�0��Sw�++lUR�P��������y�8�也��3�OR��������#s���3Q�������{�@���k�'�P������l:b�����D�����;%�jt��hU�I���f��n�ܩy����ק]�@������`�7��uAvx򿅘��?�~��Ձ��'��Tpj�(k'Op��5���O_�Ji���J�Ď��[���Ox~���UN?���ߦڸM/͈�����J$Y��Z"pT��ڠ�h��ݺf����4Ӭ��P�9W/]�ʥy���#���\~�|�Y=� �/~��.+�����[��zm��f�ɉ�y����}
�H��r���wಌ�C�s��s<�ܓI��>�{����?�j{'85*�G�m�Xolc-����f�ʜjbM�k�4I�q9�jF��QDܡv~L�Q�㽥.�SY�(J���Cf�f�7��fW/�cERT��~�c~���_��(G9~Pr����o\c5�э��d�o\����GcD�	���A��Y�������X%��bW8��/���	���O��/�s�"I{)���̟������_�wq���1΅��q���D���$�u��"/U����CIO���c\ZҵUN?|���2��G���ʣOr��'�xg���}>�or��[t1H�b���7���G����!�V��b�&���[����o6    IDAT��g���%|Q�)E^�!��Y[�ڕk��w�'�^��	�O�(�,���2N�Izn��\�&���\ӹ=�|��jַ�
N�3N�������ʐe�9{�i���L_#o��Ԝ����؇��*��m��i!')���ڛ>iv\g~�\��wW/��}H� 	��"C��xd�c&b���#<�cGxdK�H�DR@�$�}i�t7z_���z��f�?��R� 4�D����.�y��s�gmm��h���"ssst�]�f��� �$���+��ш<�Ɋ>.	�6q����>��1_�1�O�S�����O�y�����vST�n����J)0`]�$�����}�g�XM&�2e��j�	t?�E�������B��F�%R+T p���ɾ^3M��NCK�Ԛ�����/�DS#�`V`F=t�w,�U=Ӟt��oN�L_cƁ��N��b����z,��N���@K��ZҬ�xTRd#n������Ivnq��1�T�$��F7o��JDai�-�8C�e1 �.
��~���ީ*�S�� o�ए苸D�ݥ.}[r��}�~�� C�Li7$͈��&.V����n��<�7qKD�S����V��t7E��#LQx�H*:�9��S|���s�)��Ko~�[?�[�/��VDhy��)yE���Rzm��ຮ�A�l�n��Ggy��&ͅ���7�珂��es��r��/����@N���&�fDi$�aB��h���2+'��Zzi��$�>�E���7�ijV�0W�.�d���ٻ�Ecn�7���X:�	��ƍ���hx���sU��Ϋ^
�E�&כ8��B6��avR���_��W~�i\z�#�/mq��A��s�6�;)���������9GWk0�}�7������3�!{��<-0��DK�)�b��e���<������Ga���[̧G8����3O2��"Q^r���&o��Oll��+�XT��a���e�,:�p��\(3�ɀ0tt:rk��3>8�)�C4È60�ޠ�i�j.p틫���m�-�EM��#��pj/������ѣQ�UE��x����tD_�Y�HG�@���H�w�)dY~�	���L�wc�Z�O�gK7��au�����;}o�li��y�ߗ��]��Cn������ѣZ^��l�0���;:��~���>��;���d#�t�19aN;�8����$I�D:�^E��Z����We�����iG�d�Es�C{8YxQQ9I�z�AU����`1���D�Q[M�0�h����yxO����h'(�t��@��q�I�r K������B`%�٦|������
"@��jkY\�(��/H=�ճ*�� ��:�F jF�:73ml��P���:��v"�Q�O�&猛vh��k�P��.[XL�EU����5�/�rճ����:�ݸΣ�G�r�4[W֐��Fl�8��T���$�>�.|v�^o�Jܤ�$Qͳ�m.,ü`X(ʊ_K[�M9����x��G��c��ɥb�k/��覊��H����e�x�����4�l��p�^�"�c��;W���T>�We��t5�a��#T�g-�㧹��9��������|���\����C-��e0J�ʂ�T4u��`@�4��(D%�d���5��D9� w)��#��״v{��wy��'$���lݼ�������y���Շ��?c�)]�hkׯsY9�5�4B)DŁo��8O�#��Rzy�V��}���{o�C�Xc��Xp7��O���/q���g��V�B�p�JtP��J�׵�Hz8�֊zO�X��=iH:DD]N<�$K�K��{����`Gܙ���"��F;|������{�nң��{�Ì�n�,��KO�[��a?'O�(d�H�h�1JI�2Ñ!÷^��^�V-���[$�e����SϿL$����/I���?��~�eO\�/ECE� C���Z�O:A����ZIB
�ҙ��?Lɒ�a;�'E=�1%6�g��E֯|�f��}Ϟ�����]����������
e����C�!m�VT������(�*2߱Q�0x����8��9S�U���l:Ҝ��M�<�&X:�,�^��� ��;�\�B�ґ+��)������cօ%-KB��"�(��PE	R#��sR�ZTHE��(}Qf�$��@�h���m���yIo��g��޺�֒N�ñcG�t[t���(y�������ۻ�����8!X�4s��4#�`�2A[I!�WH���8)��baV�\��
[�*�0֢���I;�G�H�%���n�s��q:7}L��Ɛρ�����w�(v�����������_"����*ZSW�)|�5��7�O�"�E�+|���/s&; �@<�0{MϠ6{��u�\=b�
N�q����:��U���Xߎ�K9̅5�.���+���������-�l�H�4JI��¡�?G�����¡�#OR�=��C����p���&�������׹���<�����C��}�e1d����9��I����iuڬ]�����a�{�]���3�{����F��C/�}�k���K��%ҥ.�l��R��z��7�P ]���/X�-��}���U^�4Ɲ.i���5�	N��Z��|��(c��U�~��N����Pin^������Hy��<�5:����|��_����%�֔�v�����J��Q�M�ݞI�ی�O��u�����o���G�C�)]��V�� %�;�l_�εss���)�	a��P915+YQ���UM�ITu3��dE��i�Z��h�vo�g�X쒦)y�1*���pk������<��:D�!+�e�颴$YFiT��Rx�Kc��#�[jr���w����a��g�Etcο���{��L��ǎ��j�c��͗�8_(��5H�0�(M���������~�=����f�F�$}�>���_����I�}��<��1����b��O��"�%&�R4�+� P� I Z�*=8{oBH�*�w��B���^��A�3鴩��i�K�����Y/W�$8�(�h�5LP剳1>Ǹ�yB���� �>Z�Řɮ�l��0fBe�$	E����í[7i�b���8�z��N�v����<G�e����ǰ����!�VU��;�L%�X��>p�i�	V;	����H=f:�����k� �!�3����=;1�m_�*O4��'������+�@%T��A�@4#���I��r(��y�B�J�N�����D�8�����m��y���ń{z:bE��@��\"�"����������4W���p����y�4�>��s�d�=t1R�x���oc���ϵ�s�S>��O��	(GI�H����Ƒ����z��瀡�]�pī��?��q���Oh���V̹������s��~�#�Mn���O����9њ�W&��c�y_�SG'������F��
=�.�M��}�ֆ)NG�EmNe�	�7ЙAE1�n@+��˗�՝۬�.0LF��1�pPR�g� �_Ͳ�OU�N�$H���7x������R&��=��MZ6g������d*�ܾC7/�E5�B�q���t�K9)v��0P������W��3O=F�F���s��!�����m6vw�';�#��}{�d�S��&Z5*��	�
h9��*�b\�� ��XIo�can� 
���b0�y=u�* �1�<gX:L@���IQ+�C��	if�����&;*�dA�����C���~�g��E��C66n�5�~�K��0��S�dyBZDbB����O��"����J�4�� d��Q���[��<	5�M��a�{�lc�V���sr��G|��y(((L���
����!���Eum#�8ms��_"���d�Ljzf�M�����{=9f�ă߯����T�f�?U��3�BV\�|��A���s�$G�?�<�RQ�Jt(C_H�h���~�?�o��Z^Y�������{�{�a��|�cǎ1�����G�N�$�ᐹ�ZJ���I��+U+�Nr�J	�RH�q��﷫��V_a�5���z�:��=�3�L�������??}��X�$����tE��1���C�W������v}��f8ʨ�8x���T^��1�@�,z����wE���xǹ�/�'�6����Ы/̨�´y���ل���x�~�>[!e����o����I�m࢈���\+-�~�����WA��bSR
��$��i!*��:ΐr�&��Rw8��	���ؕ���˭�]:��������f;�"�s>�-�7wnnp��9"�����X��a��M�ݸo-T�P��� S��:���u.�o��V�f	�N��'%т�Q� ���F�Ҏh�HJ�S����P��� -|J�{BL�';lap�ߌ[�����`��,�癋�5b�C�M�n��C�EA.d��^�H	_�(�Ƥ�ˎǨ�_�՛gLJԚ�o|��>���.��'\��,e ����7H������7����3|���y6v(�׮R��
S�71�B<<�G(���M��>Q�h6�)���e,.w(s�����g��-���o\�d��#� $�q�Y�(1N�U�-+�D�C
�2�Z
t���;ذ���2��6Y�I�ls���o]�S�������Cv���]ύ�6^ˤ���ˮ���	�8H�?�C�WWi
ɥ��坟�-�AJV
:�>�w����|d�߸Λ�7����v��~�g-����@q�u�RW�O`�d��*�|�Ez�\!$j|�r��$��}n�����^9޽IۊV
|�u$�8:B����
l1E�cU�����������j����o��R��O��E	G�;@i-�`�p8ds{�f�I�w���]/~#{{{�F�G���c�`d�W��T0:=�ui�W�z&rw n�������~��dx��/������I=���>�q+��2!�M��
JT�eI@�K���E|��uΓ�j��ɧ<ۃ��{D_q����Si�{u+X�x�O<�/qPꟺ����ߝ~�jQ������V�čyvnor����(֨f�*@G�	�? ��#�����ѐ��Q�Q�O�s0�j�]%�;�&��߁��F;`��ȵ��#�r湯3�F��C/|���6���/�<�v�'���o�����vv�������];���=�
��q��8B͘4-y�������C�����	sI���$B��7dny�8Rt�}z}Bx��DZG�Z��ЪM@G���� H�zX0�6J͠,:M.'6�Q�HG${CzIJca���p}}��lD��DQd>5QGf� �htK���c�_�4^'A$��ǏG�������-�;{ע_����!X�F�HF��2��"�7�ZG��G)��K&�2�8�:����;S�б�7�3\��ӏ!�H6�(��,�(E{�0�G��n� _��r3$�!y	�$'��u^�p� 
/�,Z�V�P9B-}AԠ�\�!�
�e��'X�=�O=�B����wQ�G�x����#A�
��w�����[�#Ca���#��K�ѥ����[4Q�Q���e�ʲ������w?e��yYŰ,HZݤ��a�>Ri_u.@*�FW0�w����M��r�@_�#�d��ʘ�D}�1�M�zw� ��g��;]1 �ph�T�a�(i�4����Ϡ����
��������X�ہ��P��S�[_�O��=)�2'�st�X^^�8=�"���i�a��ш1E���.�v�SE��a�!�
6Ձ���5���)�e]�>���B(_nܦ#t;c�k���>�����������E�W�EQ U@�lќ�%$)�,	-��{D�����������]��U�����Ǧ�y����9=�<�1/Ϝo��_�<�q�痤�H�q�K��cy@OğO�^�x��~đ���z�㲂�����W����\��ٟ����P��p8$3PZ��>�"��z��g����9�,�pPCd�C�h����^b�����O��G"���D������Ar�Cn��&B��\�9���ȩu�8��^)�
4^Hb�[���?�5���3���=��ӏ�&\^�Z�6I�:�w�CG!&�y�R+�/�4���<4��G��� �0ړ�h)0*`���X8~�k�?a����R���䍜�Q�`}�ha����$�h����#U�3<��"BH\M43�>��檴@ۂbw�a��d�����%kJ�X���3Mn2�#K݈h0$
C�V��x�ӝ�cA+�Á�ug�T�R�8O���s|��^��񭗿G�m�ch����]�A�������}��.��%����<#��%���^*�F1�D!�@I�D�$4�ڔ���_��l�X}�I���<����~µ��8y�$/��-�VW�]�@�v���8WLRG�U�)k��bV3h'q����PЌ0͐AV0R��6)G�E���}�w_�K��kF��>I���Жt(H�WGl(E�,����>�V���>n�*UAn0x�/g��]�]����W���!Bz�9���������"A����K)�	��,>&q��nݕT;A�����s�b�wʃ ��nG!�DA�(��WQ���L�em]i���G8g�Z�:]���۷[YK�*�W��v�N9;���3�_1=�= �1��W�^g�g }��L��N0�M�L}!%_f:�&�$�H�z��|��ѐQ�������!'�p��tt���W9 ~C����F��9����H��{�o�A��ѱBx(�X����� t8���>�FLZ��9���Y}��F�m$Y�ShA8��|���<���oY����V��` A�R��nϨh1�w�X���.�`m0�ї~��/~���<z��+_�%�}��}�љ	��������ߤ@�p�H87K<1����F\�_h�������/�o�៰�����K,��G��"'���bg��)Μ�u�����$w�h�Xc)�!��Ҭ�/���GEh��(>��9)�"�_
N���;4�g�R1�0s]N�s��-��=�>�g��0�׾���;؝MO�,Ę�n��`N��`��[��HA�|�Q�q��Y�~���c�������>�l6�Ɛ6%�@0��Dq�0�@��AUu4A�����y��6;?ӌ�Ä<ω�o�-��w���O��%;f���;�/.0���i�cG	7/}�ƭ+������-�tDs�If|$��%v����Y�:��(Bz� P(i���Ď�t���v������/���_&n���O~�ګ�s��y�{�a6�����ˬ}�k���)N�$�#����0%��h�tBD!A�k�G�-s�o���=��@�7@�9�=��|���/(�c��$؆�_����f�`F9���.,��S�ٌI��4bhMU�:]�<�k����O_�ڼ�Cp�����C���]�l�#�VR�eQ�&����8TJ�%nk��{ٽ�/L9�k����V�8vw����A��vU�+~�%�)O)_��9���  P��u��,��YJ

�<GBGcq��fF�p��:f�4�y�#f����U�����M�i?#�;v�X�\i�JaÐ��{;�lm@�0�i@v�:��}�A�3��?S�:��9���jC`<�8���?x�i�t�u�����t�~3�2ԕ���5ݯ7&ο��V_s�å�~�p��Q���#6Ҵ�+,�Y��w^b$�槌�7�4[���_�%���b˻Q 7Nf��E
FV����ϝ��_�3��}�r�F��{|��G��L��w������T��]����y��.����W��I�	5��f��Ch�峷?��_~L��IT4O2�\��S���#����?p�S�}������:a��v���y�*777�#�YXZDJ���&K=�(%Y:�l��<bi��O�XX�r����Ӈi��x�}��]QP�YWV:���n���S�B-�9�۫^:���th%P���!�(X�|�g����Gx�B��i�B:�"�
�G���A��	�����װwv���#?YF{JҬ(���e}s����i�Z��z�Cc�� Ҁ(��
�7.��O�q����)��Yh��=Za�C���&Y�&	�QJaJ�eQ �P{#[KHk�x��    IDAT)�Z!(�P�l:6w�������o�0֮���}��@q������A��}�����d�Ts�!�nV���{����vز$Id�e�d�cGO�H�aF7)%(����s��	Ոs���o���r�:aH���YZ�y���KYN�vsӠ��UQ�NC��=ʍ��1 '@ؿ��Ի2]��e��x������6���N�V��H�c��s�R�� ����w�^窟g� ���5U���o6��y>>�p8dkk��r\}�GI�h"���n��b���gq��,s���0bn�à7�EvL������U�E�ϒ!���Z9�B�ީz���� /���RZ5���:
��RL�;�~�)o��I4��z����@:�5vlt��JY{�8'3�Vc��ţ!h��	\�4)��>��=\VPV��F��cdsB'Q2e��J�@�
��ö�s�(�������<����VW6�C�PCd�bg��% k�1�$*jS�	BT��[K�A���-[��C!Q3����:���"����ϗX��t
��>x��>|[:V9I�`���Gy����Ïq����I�����w�0G@N�EU�E*QU:�^f�w�R^�FTyj����K:+���P{l|�!��g<��\�H���$�<�^l�]��?�s�.�eQ��xe��Pѿ�5寝�����%T����E���Qڋ]ַ/q��ߐ]����~�Nc��T|��|�W�.�O��{�P�H"Q4�aX�n���a��~o� ���ńHr�p��P؀���v��v�Ao���h6{tv���s|��΀�_x�G���7��PC"<��ŧR���J�s^�C\�NE�(mP�C)�9i Q���?�W�{�	Z�>�"Y��\n�҈�i�4	��/����7�]M�M�LR�LP��̯,��l3�ߣlǴ�g ���,	U@a-2�#v�ٕ���p��SdW�����ϱ�?{��<Iwa�C�v�.p�����Y��aR`e��y,ZJ�0��1K#�y"� �ΐ�
B��d7Oy�_��:z�=#h�/�g��|��zC\�!#W�� �r��ϮF>O�(���	!��� h��̯�D�*V�[[��-�p�,�i�;��HG}�ؑ7���\�$N���S�!�=�,A���g��9��=J9zv�S���_�SClC�1���-*Ii-��� SukX*��^�/*411�㨿r��L�i�:�/���o�@*DE^��9
��]�~	72��eH�֖�r���AE����Y���dC��X�#�<O)��("Ԕ��V��Bz�^��}C	(�,Kp�H�e	iR dD@��%+�j��0�z1A �Ԅ�!IS:�s,./���0f��Ė%ySP$C�+"G�;9��(+�x=�S�b<u�C��B^aP5%�C8T��~vk#5)"3S�3�66�A����q�m����=�v�l�(R�7Tz���d�ߧ�SKʴ��$�F��xy@+6��
���w:4��qYAosm� A�
��¾�=�F�Q���Z�I- ^�`<��@;����]�U(IEw��cƻ�~�ʊ��R�ѯ *'���)$RP�E�4sq��g_�z�S,4x��'�/_�������@�ʉy���i��{�"�;�ʢ��cG���27�}��sW�aL�q������
�B�nŤ&��u�����N�,�>u5�x��C�C`-E�OC������o6QY���˘�5\�mob�!I���p�L��=�+P�8k�)B�)u �,GY(󂺘�9G������	s�{��훘�7���l��q.�I6�q}'�����cl��݂�օ�7X��}��&)*�NBas���ns���|��|�����tV���r��R����Đ{n�d��Om�a~1�b��{�A��������4z;���(�����}\E5j�2�2��1U��r���}���K����s�,�8����S��d@|��C>�[��-#�T��;�cۂ�����a����,���:�;1�?p���*ݕ�X'�F�I��R����Қ���)��o���O?#pz���q�3��*�� `!Ɣ�������;v�h bO�R$�o��0�h7���ns��T����ǚկ?I��������VX�a]�q*�sY�����b��,5\�fǽ�w%'czt��4��Z#]��a<�ÐB��°�$�A��1�L��\�*fPQ�AP斲�rT)��y1FZ�HS��[A R���*ٕ�BIN�8����(7n��ڍ���<��󤫤�u���t�qT�
��.y�Q�Y��)q�t��k-�����e��|Nװ��������Fu��Uw��g�j#?>�Os�C�f-f����$x80/-����>�����U�iP�kKJ<���q���5�t��>E�����b ����
�{�F��:=�~��{f��J�E�s�1#�ϑ�(�1A4����B6Q�uT:�����g|������~;�)�@�12D�9��hF�(��!�{C�+O�fƚx��4�1� ����D�w� ��g��-���DG�0*i�P���`���tH$��S��P�DYc(�A
�{�k��i��~�PHr��V�%�<�\�!�e��5�����b����e�-r��!dC�"�!��JJ��I�(-�"�)KK�����P��F@�rZM��?`��͝뗘�
D���Rn���V�����~@o�g�*��OT�޶2�Nz�Q8�Rh�@iA J{���ܨ	��t@�!:ܥlj�nD�u�K7>��:dBPj��a�8Mi4cF6�9��~�oY>q��>�����U������1�0�`w��J���	*ʌB�+<��o�r�wn����ߢ��Ë��3'���O��W��&���r��r���$J�1�_�@	��EK��;@ʋ_e�$͍���R>��k|��7P�.sǎ�ͳ��S��'O�����ǉ�\:���A�ocsU}Ƚ޿��OR�Z�%� ��}���C�����wYZ�V�^��IҼ������V� O
dn(���d��B�bW ������U���hx���A��9��H)��wC�����8a���X�d@j����sz�P��F��&�ҿCń�A�ٴ�/j+��u�UW�K�d������R�A��ڎ?ƉӧXZ�C8�v�Ƒ%)T�xBͦ	�( �b�"#�"�2'MS�9����RE�U�S)k��X�E���ٮB{} 8�&�Aܤ0T�/(ϞV}q��:��y߲�8b��1�#��I�8���줋/5�5�K}X �@i�8@��,%�n�MlZ�mm ��{V`�@E���"�O���S��^�
A���������"���wS��/)H��*~�]
����	�IA�� HO���PVFz
s�ꉞ�4��2瓵�ӓ^rX(oh���Z�vb	�(�fdFN�YZK�x�G���g.���׹���,ʐ8��+�I�Q��g��0���A��sE�4��N��ߟ�����!�Da���}��y������|���&�J�ʚa�t�	��{�+D�:��,l}y�4����:�x��Ͽ�C�}�@�(��� �bYz�A��1�(Q@a	�	<�ve��/�r�������)J�1���+\�����c,�lw�N 9|�Y�#3��F���+kp�ס���C^�<ze}d���A@:%F�h�qJ�m�X|������=s����A��@��@�$��T�������?��� ;�������<O�I��~x����XN�w�f����:Y��)Z)�0�70t�� �ܼõw���-��佄�}��7^����d�($��4�eEXSm�JB����[DNn2��(�Iɨ�HҒ���֡�,��7��\���_Dv�<���9��)�E����w��¯���k�Xh���"��F\9YbR-�_*�ᐂ��<��.ŭM��\��]Af���c_yDb��1�eH|�0�H���Cñ4)��5p�d��ewo�������vC*IPQ�K;ٳ��z߯w�{��L�7�t���[�~���*")BJ�2g/�Aff�<P��P�u�8�PL���)��D�fզ�lL$��s�U�EQ�1�,-,�qg��`�RR����@��O!k]�^?!�cʲd���
�Q�P�-���ʣ.
(�\ �&�c:z���3�^���˽���@����`�'ol�}w��Ӭ>��5�A5�`���Փ0�F�(��݈��wq;%�A��,��(���|���LI��c[�d���K�}N�Hs\�\�T�i�FPk�:O�0�j�r=h�'��^�A��f�$�S�,��B�de��GN�ԦQ
x�9W�����:%��A� 8�#�4���j|_�8���������o
�� (J�vL��1ZaL�����~�:Q����j���!U�h�tH��P��d�N0J�n\���ϱxh�~@��t�VV�ZXD�!�R���e�{��cm�-L1빹��UZQ8������u�e�E^��Pj��� \���z����9���5�^�@8l�"c4HhG]�,�ֹ���ހ��@�6C)	*Y̲,�4����`Q���Aoș�����߱��;ۜY\FHU�F��-K�ސ��l��6��ɨ��_VYuj`,����0�Zh����"1��(-�]�����=�����m6��`��E����:n�5�&���y�"۾ƻ?���^�c���l\c���`0�Y#FROֵ��qH�hJ�:Csq��� ��t��˔�ZZ
�I��`�!c0iF#��~��/
Q�=mj5�ZH�ҞpŔdiA^��Na�F��j7<#e������K/q�kϣ���sor��7�����יo����ׁ�)$�>d��W�"֕H�kZJ)9|�qμ�-�����_?�Q���%e	"1�hd<�헉�K׉�P�e�!��F������=�C���@��X�ua|0��g}��ViÃmtUE'u�8�;R���=gz�6����p�����Ya��짾�N�9J�����hi�XL^x�nj��BNݸ�~|�¿�����Z��Z���&7��"Kr�~q���n:�i�ۨ(����@���0��k�B|�,��"�Ch/���/� Bk��V*O�%=u�qvL�%���p>-�e�����(]�O�{Ů�҇�c�~�8x�ZFLj��:�=���A<�&�����y�b0��D�"�P�\9�Q��Y�ՑI�$%��Yx2�Pi_�dథ!u)Y9&���bń�WX����P�U=��>�<R��08PU.�"'�F���4��p���J��(��i����S���tF��urI���n�tL(MBD# �����O���"���gt�A9C�ea�/֬ #!�yU�3��4Ŧ��!8��_����vi/����ɉ��ԩc���D����mFWnRd�@��!��*GWX�i��%��DT��Ջ�F�F��c�y���u�x�UT3���}�fѥ�a�d�Hpti�ls�s��o��oн�P(-�e��[	�Ä�К1���NQM,��|?����MGN��N٦Hs�\�Lی�oF��{�Y�q%��(��1�QT�3/V�|1��X͔1e}Q�Px�1���s�I�������b����]֊�w^�5�O�$s�C4҂��u������8��.a�υ7~��R�EL4p�oޢ�dE���߸�j����:��\�5�����aV�8���nLjv�!���|�E�V,�7	;]\����0R4� ��3�%���B(� )H���!H�9^*(�lؒ}�3w�i�<��<�$G}�^������_�������ե9��A���I����A���D���Q�����x�=���+�)Cd F8k(R�f�uO=�^X�3J)���utY�m69.�^`ws��#�PV���A��DJ�(xbg-Ri&�cwG����ei�z���;w�=�w�C
������9�ܒ���Le1�*V�m:��Y\�S��Lr5K�+o3��Σ:j�a��TdB��QD�s�ܔ�Β�G|���t�-��>��t:s���W�Oun)��:���cq�;��X�<G�A&v�9O2f��8��Eh��U�=�&f5�gBK�&�`Q���PW-�ιWE������^kb��{C�f����먿8��67)z�~B��a@I�$Ŗ��EVkB%�e����%u%ҁ�Uu���*�d�ԽY&�4�:������c�>'T��n��!�luj���0S��d
)}�ԥ�gy�^J���|����%,���y�/��]�QiQVҍ���HK�Z��p�}�A�����!a�AZ9W>�Q<S���Ĥ�r�_���9I�i�!��9w���8iK�(h���fȮ��F���H�a˂n�"��P�\#B�r�_5�!����$�Ԟ{?+�o�B�m�)�#O%iKHo]���/���[�E�IM����Q���&���>%p�;��y^k-�X��D8BL6���`�2��u������?��s�*��}���{��{��w��C��:�ɲ���h̏�����0��5AQ!(����%e�V���h��B�K�6�����̙�<��C|��C�����d�y��;�]b��ڗ^�n�M�=��(	�4c�g�x ���_��1�؆0I0,SC���)��{wumY�K,w9�?��YE�p �U]�q�ƽ���>�[�7�I�+���w����}@�
�M�]j���������+\.a7Ni����c>���Y̖���xᥗ����%�v�y�U$��c���ů����T�����7�b�*d�H�V �\�fI[Rx����R8K!9�Pĺa4�坻|������`�p���w�_>��� f�}%OW'��9j�����5����fqSJ\��TUܗ����C���7�����맧�X����y��l:���Gf�pX[6�O�1uӖ@n=��3mZ��A���X�9�yw�G��P�uk�e��gm��̌��x�2M$�C�|ȸ��Td�cU�Jk�RZ�Y��C$�R`?�(���r����N^�Rb��R�et�5k�>*E!9:8<�29P
|����v�B�}Du��<TR�"�b�N�j˦�.|1FB,����gL�:Y�
�]1����J#C'H�b��� ]�l.�������/6�r�<ӐK�7�y~6�{�_<����6M9����o�a�EfIT
�!'�����L���<�2c�,�+r�V����3���\���:�-��_�\�ÅP\Ô$�P*�\:���_���ܟ߉�ô��w�D���]�E�xz�����5O�����F�;���V\13FV�UƏ=�%RE��,�,�nV,q�Q�k��/d�����9)�����T	�W51�؅a�,~,f�JK��&�G�ؑOG�A�Lnk'��S��z�r&�Kâ1�T�%��oa��.Nn�H>�o&�TP	@��CV|J21n��������R0�j�@,1�)"�A	�КJ+�wϜ��EG �,f3������G�+W���O�ܗ_`���~����x�*U�%	OGbX��0
/�nv�V)e��k����!�K��я#Y�|n�%i�o�+��Jvx�����1���8�!ƄI��Y!�d.F%���+��ft�1
A������{n+�������7>�y����v�/�5������pcvċ/����1��������lD_�AH�Mj��I%�Q+��5����Gb��>!�P6�p"bo��o��}�3�p�YT|����ջ_������{?�?��o�����_Y��k\��ʒ����2!51Io�­{V�y��.��j��g(��z�/^����#֫V���;N~�6s�p��W��mj��W�� ��o#e)� O��T{N;/������7��b����|�C$A���N�#k���F+I
m$meY65���#r]
'�Q��J�����rb�[K�H�b�6��7[�KS�g�T�'Wb�S�a�MM�q�����C�9�8��1�X,����HO�2*݀B����^)�҄�BB�֍LN�,+    IDATʰR�ĉK7=�6�,�����$R�$3p��l�J���Q�"�B,"er�-qz*
�b�"e�C*c�L&R�DC��X��j9�N%k�Q��c-K�s��4#Q%г�(D�X(���cL���`E���#�h�0��Q�؝B*p.@
�ō#9E*������l��.3��X�Jw�.f�Y�<�\*8u~�&�%�rulWg�Z���P<������t1�Dh]`�I�!�(�O�ЂK�o,o��r���"�,%��(?ga(	���Y��LD��J��{̉чB.K�(�dQ�u5-$1F���$C,$D(]�3Z�Z�	1L1���S+��0�:��g�b$�@d$YMp[=3%�<�x��{�P����#}��)9*�6R�R$E�h$"%t΄�Ok^�^�Ad���n5c�3R��+C���G�i�&9_]W
 &�lJ��#;�
��L�@�@{��Yp�kj-8F:�Q��	2�h-���RD�TF`�BQ�d�.�a�Xo:���!8L��jV4�n��7��������;�����>$��Ȑ3i�3wpS6�I�Х�����A+�����!9r򄍣2!5Yj�8rm�Y��������U^��WpY���w��/����
�a��?��o�#?�������s6���2G�\�cʘ��9]o	!��FdA��3�T�F#SFY�].�]��1
9-�����R�j͓��3n�����ǚ�&D,�'J��I*��Ժt�OU&`X^��Z�d9p?%�~�?|�o��_�n�y��3���s����&$������G����)�޸���)o�����*<|z��/~2r���V Q��U�݆��^�w��F�R���;�,z)ws�I��<O�?q!�FY�@.&����&֛-�IJ-��$Q:�"s�R��*\�W�T/�B�r&dMkZD?���M��K#q!�B٪dM 
whV�Sɟׅ߮�a[Ԕ�Bu�j*|���`1!ˁ��ݴ�
k,�H6��z{��5M�$0M!(Ŀ)I�*�F����Y���舗y����	�P !���R2����dQ�{�[tM��iUJB$���)���@�	k+\��}��iK�<�`�+��B!�%�(39��4U*B	��)�(3w4}@&iA���8R�3m�e�Ѵ���k�y ��S Cq�۱@��Ib�4�&�Lӄ"	l?b�' �0m������<��\.!��J9���\�/-.HqR�ٱP��|��ՊN�Z��Fƀ�-5"�H�i�1Ő%�a��c%Z@�)$:��Ie�A�c�����D��Y��2��X$&KH��}�N�DSѧ����ƴtkE�(4Y#���3�,	1���$&��8���H�R���e���� �����J�V�����1��F+����RItdH}`;�C���ؘ03AkB@�"IC��twuŘH��z��̀-9b�CJ)�����R���E1��%�-O�a{��Ϡd;$��t�|n���7y��^��ɚ�=��T)�>_��]�R�V FX�+,ݺ�X5��0� (y�_ 
)%�:�g��u��+����>�_�"O�f�k��|���TY����w���h��;�q�o���D�܍�\B�|v�}���E���e�zX*���g<x��������5!Ó�3������8��[o�@��A;c���Z��QX�J[�q�ږ���z�iR1��#�莟�Ο��?�9XK;�}�����,�!н�!/�� �贗FM����V���ȹ2Twn��K�����'|���{�x������撧�=�z乥j<~���a5������v6�9�4?�?]qs~�A����w��q�
���C���d�*��Y��hu�B=���Q��?���B��$&_�_R�P�.f�$Yu�.��'J*�12sPW��	B�l�6Iκ-���b���!tם�qrS�]|�e� ���4o���a���B��Q\p���S�0⢘��^�ۦi�r���~���w�y����Ѷ-z�ïU͎�|�K)"o�6z�-�v�ߤh�j����B�¤"d��0�r���Y�:"����iIƑ�%��#��0A�)k�X:�=\2�ݦ��IY"�-�k)H���l5�(��JwJ��G������!9[}Z��9�P$�l���iC93�.����X�]z��)�T"���<�y�����r�Τ��&�k�K���d�"��OJ�ֈ$��c ň�g[ӏ1GF��"#� "IfP����)�C D_�T��4�'�x�5+��� 1�&e�J�
q��'���B����@���U�D�&���E�\�ݔ,�H�Ӏ�j?#T��QΤ�	>��3���*������@&O�T!�d�l�
?c̎U?�t� jŬ��ĎʔB��Rrf�	�)��M�v,d$i2����6Ƒ��h�`���*�6��(����+Z֜T�����5��D2�݌��Q���r�o���s����a�Eݹ�o�@�-}��-u#�>�����w��g�*%�� �VȢɎ�at8W�7Z�b�{���/�̗��:��!=�_����U:��D�g���D�������Ot?����+���0hm�1�c@�Dm��|Q�.����j���1C���@5��]G<M�`(ZfQ�\?:d�=F��(
�zt�U爱��r��_2�k-�mW<�ɏ���c��3�0�u�ȴ�$-Aeb���F��ظP�Q;���w����s�^��w�w_��u�����{\'���p���e�(ҵ/FN>`��k��{os��S��!0;\��5ܚY6ܾu������ ��㆖x�s6�1on~��"��Ŕ��g��x�c���+�����EW��������a�.�.r�{|R��&��w���,mME��DE���s�:�b	.."����`�]�/ͯ/�B\~�6�ݿ�^7Ʋ�H�+$:)UY3��FXirY���pyDƃ]Y���#�r�LR9!vc�B ��r��/L�'����$E��Q�~]��"!�HXk,�jB#�����ad�>�'!e�i�p��QMU� �rp!N�6ʅ��Bb5��1:Gm%�*3���H�@MUzv�4�mΊ�p�E�#!eJђ3y�̈́d'�(���}�0�֠2Xa�DM��d���!E�CT;G�#"���)�l�K(t.@J��]�w5A���qt@�6�$��s��9<Zr��N�7�i3-֌JJL;é6g��(�0B�e�0�%Y�)� �w�q$	m,��"���l��ӵ�L���i��0�Heĥ�$**S����d��C��552�s(!�m5Y'VcI���V,[��l�Gf��9bU�w %J)�S��ԍa�
�R$��&u�T8	A+R�H�0HEv$���i3���O�1�����/��UVX;��r�(K	>�����!� ����9�/q�������>�s;������"�#m���H����?&��ES�����h����pB|ʄ�
�I������
Fǣ����7s�}�u̬��ZTS�$$A��[�køb��C�.=c����*D'���T�PTZPk�׊m�V��g�(-88��\A��%�����B
�uU�ʔ�bB�;O?�1�6�=	���A9g6
tH�9lʼ5��UE�qB�ʚ�bm��*ֱ8#���1�;Fe���h_h���ȏOm��,k�,�b
�^�9=a���Wy��U��9�ɊP+�چ�T�zɲ�����Cf����B��ß3��U�z?r��M���Y����I)?�:}�h��f������r)���g)�(8��K�{�im�����$ŕFshC�*͙����랡ZpX7�	]SU�Ǜ�Sc'��}���ra�SqĤ���䫪8ؕ�gI��k��jG�fUU)�P���#;T�|�����\=:�s��'�KN�/P���wW$��D��������_6��+E��B��$^�=O�S��54����$��=>��t�*H��~'-���9�=��%�4%L)��R��d!I9��7��B��t-
\��FP�%&$R߳uO�Y�'��L5m�i��KF)�,?��r�t6&H9�Șv�y���f���.�ː����Eۮ�.�߬Jk*�A��rNE�#1l-qc ��( J���kܸu�7n�9ߒ�Sw]��t�(��6�K
;k���� �,�C'#����4 D.�gJB�|�~
RH$B.L�������q��PC$�}����d��h1�ms&�ȿ��L�:����>1�7,�Ī�q�F���i,Ѯ��_��2N{GҒ�G�5-7ma�Z_����Aj��֢�Gb�Xk/ �1�黛�9G������l1g��t]G����1�|�G���i�3�c�$mPB�住����r��X ��;�Œx�XՄ(qkǙL�9�>ꩣ�+���I��EI��!�;?9�	�4����99�������ӿ�O����Bl����	j���R� 5M�I#��	r�FTG�@��y�t���rH)h*�5%"���3�J8M�D9Q�B���(3��
�ue���G��U�d�)f+�H?f����1�����Iu5#��$"q*���@j��auE�d)޳�dm86,�9��ҁQf�M�R�[�֌f�qC<?es�Ó�Q�S��s;�ɒ#٢r����/��i��`I�4(:��� g���F�Rs��-���:7p�s���Y1] K�Q�	��Tߝ����sųd�39�-Z2�I�񙭃m]�dc����G�:�����H�=�}`��-�aZ�;�B��n=U6zb�_�/[c�못P������ϸv�MӔ�����~�(�u�_OUUM�
� <�)k�r�`ִ�����1�ْ�þALb�#T��|hU�K�=u���R)ĆM�"�y3#V5J%Dn��)C4�b��^m��'F�/�8]1\T[1F�tTA��V
���|�sl�-1�@�VJr�I	lm��n�8F"��uJAul��Y��t�K6h��FԚ!�bèT���q��ΰFJ��^��QP��2�9�r�,! ��o��yKʸp3�2��,��3�v�u���cNO?E�@%�� Lq�ZH{��,��֨T*�S�;��	��(G���4�P�!oe�j���v<+Y
̔g��q�͍ �d�:�ڵk��P�jj��5�s1��l6���72E�"���"/�Q���s�޹�ʂͣGD�P7�c�d�� 6mN�bq2:²�.�ē3�_�EB��;�'��`̑ӳ5#����ɔ��R�K�.7����k�!1m�RQ������RbM�kH)��
I�g}`�(�pU޿��~��p`�or�:V�S\gT�����t����b9�p��/ŉ48��HH�81���r�w9L�RND�T� �����kt���s�{��,2&g�C�p9�t�y�mUII
��V�̍Q�u������� 2$���vל*c�JMHKd6�h�A�T��ڶ؇��gt��'��=�e=xYH��9g�X>��"A�T�XP$D(ֵ��!H�ڴ�n,�U�.�k�9G����)�
%�ZAآE�X�r�!�O�+A�`���YC�$�8��Q`{�L��,T�D���3kg*3��b�0[.����s$/H�����.V�=�jw>��Iw��gI��T�_z�3�r�����1r�kC(^fʋo�����k�4t�1�mE��X�<e�G����&	�s����½�t]�8��D��X���=}�G|JS�[�5km����,�m[n߾͛��oQi��Dh.�E{Bد!������q%�秤hj���yy>;kd��]*�C�/�/`�]g��H�.mq�!�27��«;xz����Uڗ_��7��_A�	�@$ -E2�\B �R5�.�a�%��3E��#���ZT�1�����Y���T��ҚU��w�����b�]aMN��>z��,X�MS�pJ��� 
.�]w�I���BT�0n`�$M�N1 7D�/̀�V	f�|G&AV�v#���r��7����l�,�3�4�����خ;�����;E�#9E�H��0Rq��)n zȁ!x���W%6�����Q��w��Z�ιj$Q��^dd]��'O=N�����y��I�Њ�V(=E~�r㮤d;����gl����Gв�N]w�V�6=�T,>�
/��7��_Ɵ������c^������Mݿχ?�'�|�ELܹq��醃/�ʵ;w8}��O�G�4��Ј	��}`��{bdI^H�vs�]�=�q�%��Md���'!�X����\���1I�s:���զ��#s[#���mB���m%�<E��Q����cR����H&��R����.���8�M~�,�i��N�B
�FI*�ʼy�����HzguZ��G/���p����D6�(Q:�:+Ѧ̋��8��H̉,�d�H)�c,$:����
I�V[B����R�#���SĥL�˽��ĥ����ج`'�M�!�DX	"�ܚ)�%���b($ڔ	�����S����I�>B����hd�0R�Ǟ�w�2AV��!�J$0ɼj0�19�K�uG?th�WB�]���}��n\���
�GO���͝�(9���r�	Ռ�U]B7�=��r1�+���M�^��w3����WB2���V.��H���0Ҙ̕�%�3��nq]h�T8�C�O	i+�1E������n�a����n�'i�L�XxMJ���i̴I۩h6����	Z*�nSb��!N�2�w��wE)���am��ӳ�Qԕ���1�M�V5~�elx�����\鹱�xv��x|�� L�)R�r� ��V�n���^��W��=�Ijd��"BLH�Ѧ�	Η=nGR(Z�#�c��緖�����g�>Ĉ���|��o���_cn��d�E��ҙ��1�Ƒ0�N%�.��N)ML�¢,6�%�n�o���6�U���O��o������H֗�C�4���
�̇�\��wZ�b�CU��P�#N�]��)Y���o�&��~�=<����]n��7Xg�uCV��T:ʄ0kkH�quL�0v��ʆ���*��'lWk*��)s��	9�~�|���[%�1K�rFu�:/�E�:��Wzr{J)�=�����y�>��:�Y�l6��l7=OOO�x5��79::�]�hD�4���ܻw�`Ŧ8��K��G��;�+���5_�r��G����~���SGWy���w��m�������(C]K$�a[e��9�:�>�Aj��`0�&�Qd�Z\�'���'eEYԔ�h[Ў��ϸv����0l��"jS�5l�rݥK����9�n�G�=w����P�b.���6G�	2��5K���ȶ�%���q��q}�H���L��KeY�{V��.��11�B�U
�Vl��3V��W�J3��_�.�6���O�X����ՠ�4/�jN҆s�(wQhlJ���
���j�KTg����Uj�VDJE�iKll%�g�41��1N&TI`��y2���Q�H!��c	���V�J�v�{�Y�5�J+r�$H	�.��uVEI3sU��>�F61zre
�d$Zj��l�������,�F�ud��k�L�B�7GR�jK�,f�n���!C,꩔��P��\8Q��w��gm�ϣP��y��w�%/͐�D���!D��l�.
�*��J'��̬ 7ҭWhӠm�j3�8l|.2�I�L��$�����:�S뤔��*��;����햜�>�&��R9_��t[>x�C����I��zOГR�B>Fb�{d 
ϣmfHi���Ɓ�����^���vI�e���cB���_*��M�	c��[dR$�A���(����z��5�rN��=~�[�:��.i+�r���RJt��9�tԪ��v�z6x�aK��)iK�]@�!�z/ٮ7��rG�sU����Ր0���B��w�+���,g��5!G�UX��T�ȍ�����,�$`C�z.���/��q��1~�X$�Fa&�$�Hm$ەG�~��K����QÀ���%����5��K<��1s� �'9F�,&E*&|�c�͐B���֫_g��װ����ػN��,��Y�Vl��.f�W��>;�`>�	{3j    IDATu=���-�ӳ�Sq���g�l|���>����i������D�(YKE��+�����zq��M8�n2���1R��d,Qk��
��9䬦>\r��po���m����7,ԂF^}�?�����|������淹�[��6���_������������[�����;��ᣏ8��� ?@�����O��ֵ��n���[��t���s�$�J�r.�-�e�e��Š@�p;�ZAJ��״�X�63=:q��;��F�9_!UF���O�1�/
���愄4�y��ggkfU�t$�b��\!�.�����ŵ��b	�ul� Aa��/��C'�E�!'i�B�D��u�0����f�P9��2 ���9�	1`?�SSr�,��4�����������Ĭ n�IJ!+���1�Q"��׆$uA�6�$�C �J��!�Dt����I����J#��䨓Eg��.%z�s�6�-]ױHg���A�|��IV�kŕ�0�9�COp�#e�!2��O�bŪ5+J��D�@3gq�$S��d��s�1t�����Ҋ6xfVё����iD�D5�|O���/Q����#3�cS d���('u���)&�q�\�v]..����/m>;�%`KH˘"[?��TJ�r($e+�Yk�>'�^�t�e���@�f||J�\Gd�P���(�J�P��$�� ":M�_	R�)����S,Ȝs�����0a�Fr̴�Ň��V(,$�@��G�ĬV*�h�G�
�M!�*�͉@��D&�h֚���Ź��@����c!渉�DBN
,+T1�J�U�����ů$%�\��v��=�2Id���F��W�7o�Cw�>���_2~���蒠��R��܀n[��+b�v�8tH]_�0�}bfk\��j��DK�=zx���	� a8�<�?�1���zA�[����*xNW��#��!"��].sDǢ�����b���u]s.&7�F��_|��撴)�H�%L�9ѐ���	����o}�7���<��}������ܞ�$�����y�Y��X-q�-"F�)��,A�c���8߮�砮���������c|_��BU��,���g+��1>����h�y"]v�1��w&��+>�tTʰ��@c$�c���1��mѪ�_�'Oy�O�8";�3[��Fr¹�����dF�LU��'��UQs�7o���|Ƽ���`I�P�V+������w燜�c^~�s�Ê��S�{�|��G�=z_������Ïx�ͯ�	ϡ�4�o����h]b*�pR���Ѥ,َYL>�J�t����k���~��W�L�Dܮ��L�� Ǳ���ٚ���Fi���P�K��՚\����HQ��s�gH���R �X��:��Ĝ�)�%��s^��wA��?�Nk/��5��ۋ���L�ϥ�^��`;��9�d�[�Q'�Ɯȹ�EW�9O���C0�e>I!i-�z�rV�&Dp>�B�I)�ρ��)RUئfk�*��2�<�[zi+��@u�T&$���Z��d��q�$���'��l�ӫ�J�7�����@����R+j�0����>
9����H��t�X�$#�d�HH����	vV!��۞8*N��9s9��#��UE�e�L�|$ň��ܘU\�tl�"E�L���Kc^q�A��_g~�z�M�]�z���j�H�

��ē�B�#�s8����i�2�hjB۔�KD�uM�z?6���ER�u�G����w	7��/����E.J��޲v�䭡�2Jc9
B��#�i��%	�8x�s�J����1[�k}G��#�)�З,zw�G.�~�µ���)�u�S|-��B����.z�(�&�p�f>Uw������ӷ�°��Ǎ��}�m,і�[Ӈ����~�1��ᦃ�(�����=�py�q�ѻs꘩��27�H��Ǭ?��1fr�X[#�l�2���,YU��+���<����CLž0zje��Zd���h [^��?��[_Ǫb�`E�BJ>y��ǿ�W���Hcd�$��+p���|�7dbX.��ڗx����ݿ�s6����o����������޻�	F��|^���0`�5���{|���t�lm�051$ڶeq�f9���W�~�JI��9�|�Ï?��V�q���V�fp#^dbؐa;��Bk���G6�|��{Ȧ���L*\$J̧�E�PU�łs�Y�@����`qȫ7op�d�$��	"�r���m8��y�2�C!�F��bk�z��w~�S���~�s��)���7��_��'��+�G�plj=J�$p#�T�R"U��#c���w^��m^��3A�Or���w/���;�g)��CrvcǑ��đ���d#�Lte���,x7�R��!�RX�����Lz�P�(��녌!�ˉ���x7�)K�\��i�ķ��ȧM{�'�K��#SC /���ʜї���؏δV�� #���1��,RNS�Qr&3uJ��W�������1��zU���l4�Wq��YY������Q1�GW�m���lV[�.���p뎏��c�ˆ���r��U�rI�,k!	�-�4�ꖁ5q,�BNs��LC-�o�|���1�(n�1�p��{Ϩ$1�x;����D�B/��䜘�Fk�.⇁Y���>�2#�J���%�VT��n�kE'4>+�������}'~	ʿ���&����30�t%q��#�1)3!�$ˍ�t.һD���H���,+C5�t��L%�d���F&�}���]8Q�q?Y��F�~��#_H�
���94��H1"rħ�)�jhꚣ�#NNNǱ��TQ[��j���r��'!!(Q#%���9sي�W���/�1����fF�NMR*)J�i�	�JU-Dhg5�L4:�֊�ʒ���'���?�I�x�a{rJ)��z�p���c�zÒ_9� :���9}��m+����v��I�y�5g�����T�B�l��s��xGGב�`��"q��;�s���4C��o7$%p��w��GO����)��jMΉ�m���9��"�|�wH͌q���7�{�X�o�.�(�_��o~��?<���ÿ瓿�?C�H�JB[ʩ��tqĈҭlG�:�\1�{��x�I�-]�S�}�����Ɨ��9�z���oNs*��v�k���ǟ�����#�*�O�Q��Я7�l�NL���!{Ҡbf<[!��<�l��G6>@�"l�I
�{���k/��/�t�������R�@{�7�2Z8�#��?���x�+�GK�\�C�*y *K☹z�*Fh�jA[-y��	��>cv�>�Φ����vRv�"_=HS\�|!-�L��c�=�$��3��1צ�,�վ{� 3 $�Kr� �JZ-d?P+�k�FE�\)$-�� wC4 8���fڕɪt���fVus@�FtTwVvE�5���>�Ͼ�L���R
ш���J��9N��#� cQ�C��
΢u�������q�h8�`�]!nd��n"<���s��Ń+Q2ڋ�څ���ĸ��eL,��v^�b N\p}��N�ݴ������b��_6���	���?h����}�2�\�ȔGnd~�zR��|tY"B�RƴI����$��z�j�s�u�P5!S����4����o���r�C��ߵ䉦�W<{�9��AIӵ�C���Y�Vŀz]��]W�4tfŝ����C�
�^c��8�����IQbV��h���1L
�?{L+��]9@%,��������G�߾� J	g�m[㼡ԊNKt>�A6��G�9����@o6*�	I���4�K�iPX��FL�¯��f3����"7�K��f�|���k|�\��=q���}�%R"h% x��X!h4>`�(��6J�Ge��������|��Q�ŘWKoL���_�
�!b�|3�B����2���x�RI�:8���^{���1O�<�����lF]UQ�#{K^I��8�5EQ@�1Q����qz�/\�����%o��s}�A��_��q�p��z^� ��zZVJ|E�R4����ѝ�ҩ���!xڮ$�*Y�N�>g��	'GG�J�导˭W^#Ï��?���O9�9��;$ݚU[c��{��g��R亟')�uגܸʯ��%�䣏9}~������ W�87T�D�1�щ����T���s�����1�
%-��0��1��3�G�޸M�!�Y�@L��C���y8?������'<�!�%��h�w&j��B8O**ҵ+�s�EJ:��Z"�������ȹz�+L��u���Erp@K:����Q*#�	*����ϗ���;��G�f3l��Y�Y6k�D�B�it�V��Re�=�TT��rB��W�s�>�Yv-]p���_��NGȤ ����x�p������������s�v���\�ݺ���D��9�+��y����YB+w��5�'Oy����_?�L�mI��EI`�����s�2��лH摒�D�mR�0�7�ظ��O�%�\~��9�P:Jl��b!�D p��"Kw3��ć�I��,�<�H@ے{�,�L�|�x�LN�>S��� 	p!����P���_f�<������yM���D�o�)8�良����l�J��ד�-�z�����]g,��t6:v
.d�҃;��u(GHP!&�)��r�Z���$N��Q�#����5u��Δ�ٌ��?��_'�D�v�6�;Au��Jlԕa�{�ns��-vG{������}�߼A�j��A+���9çG�M���}�?�-�	eȋL,>Q�F����r��������PZ��>	sk�I�s����?��K�2��g���)� ���j���!}�Ø�/��_��������H�7�7�Q�}��X!�|�nB^��Q����0��ES#eN�4ț!Bډ��:�H�TѡS��JFk���U*�:O�)�z5Mך-9/I���k�,Q I�fgg�7n %\	W988��쌧OSU]��z�$��qk" �ĸ@�6��ۘ��1��2ʴ��I!�C�o6v��\:�[��Z�n��Й�1t>@��*��f���"(E��,��DY,+��9*bXG��|H�V���,y��\�'�wVqr~�mb����#>:��_�U�r�C�^
�"�i��&�@j�>J�m#��[_!;x�jx�5'�+�F������Zd^\&��&�Q�-�<x�]�U�2?;�^W�i�c�k>������w����wX�/�[K�ȇ���������;�Ja�w����4��:�	��x�N���Y���4m�J%$J����p��78�}�����:g;���	-��:�yN|�P,w��>�<<;&�v�_��_�5k�<�G;�1{����)	AK�w2n�s�T�*�Dz�]�c����[_�ؽ��|����9��iN�,g�#EJ���m�x:f��jw���e}~FW&�V1���Q���Ԓ�t<���o����Mn�T"M��2g��k�-��b��y������⤉�(�!��a�'H��.:d�ύ��H��&.�}���Z�F_ؚ�Џb#*B@8�z\!i�a���lI�Kj��e\�;s�l@�~sF��l���:�q-4R��;�N��o���4��7�7v	�MN��MYnX��E3�/�Q���ݼ���'����g��7�@��;���v��.�ERB"c�d����q�fX�uCg<R%dRж-�R[��(� GS*~��!V'$YB�Dr���j�lv��mjX-��Rq~t��ǟs0��Vu�����)�����������Th�u�����>�D�*�Vh�1G'��+���l���>�2-',f�q�o;�4M
�rH���I2`/�`-�Z��d��)IZ���&�Eu���>lkg8����������r����?�?��X?����@tf��˗���g�>�/��C�|��`}qIw'����zƿ�D?N	�=�(������DH���K�������ڦ�PJ!]$=ot�I�`���K�����7���	Zm�sƘ~~N϶��`�e�\����Z�8�?�Ν;�?=������ӈHh���
A]x�8���u[m�R
aE��
�:����Z똴���އ^�i���9������e��!��Y�	2$�*�q�h:a�ޣZ��gOi~�#���.���06��ڞ�(t�������dq��|���bQU<y������ck��h-Awk�B�=�k�T�H�������Op�0LS��wx��	O�c��1i&�&G�g��4�u�UC�4��"��\�D��R�#�U��{?F%%iPdw���㪔ݝ���<����Bjj�L�����R��j�Z�$�$H�m֜�����\�Myp���Ag�匽vɧ���v깶��b%(��'M��L@��2͙�����6��)�����o�`�7L�u�>�H�B7*��g+K)��W��1��l!0m��zE�v,�KƋ=D�1~�.�ȳ�3fu����:*a2؋��5���Gh2��˿��ׯ�g����ԍ+�7� ������2��G��ZoC�w���8&���E����!HN	��C%q� 8�w�BA/;��Q�__�h�k���IS��-r��0_H���X	��]�t�6x�W�K�H���yߛ� tw��:�7� z�zm{�����*ba���B�9�p�f�,���b>E��_�) �����k!{���*:�O��$Z�kA�dϥptR��s4���zo})e��p�/�+7ؽq�$�<��S���݇�ՂNAe;�uC�Rvvv�C�X@Ӓ��9J4��ȳ�u2�4����N�5W�c��u���NEJW-9��C>8>�^��+%���%Uע�F�42��[�'W)I���!Zkf͐+�!�A�\��׹�����3��g�񧱋Mt��Mz���<��|�ߣo��/ �KFb�C���$J��J�К�L��,O�Yp��p)c��>>�����1NZ����m��q]�T̵���D\�ɣT4D��e���罘H63��/>O�Gn�Cq�u=Y�C�Nb�!UC�:>�JEr�G�8??���۔e��ի��Y^����;�<�I����E���g��m�5R��&�x
�������ySh�K���ͣ�e?�cDd��PY�h�ɕ+8�X�V�EFX4Py�Z|��C��a�%���{�*0���t\2ݟ�^W<�����jv����'��B��ќ�2'tgH�!����F*v$m�a�CY��\ �;n����$���Cr�C]�4����Yt��!|`<S�n988@�ğ���B���K*5cze�z~��?�#H;^�����S8m��Ss����8[u$*�Z���� *ʋ\��
MJӮq�f������hĪȮ���FS��{̳�ⷿ�M2鑢$�u�@����'<=9C.,�K��w��OO ȤC���(�3KBg�u�@*)�S�I��h���J��y�����{�'�y�s}���T��%6OH�� |Բv�Qâd�q���љ���d��J9�|�w�O��)�[S�Y���1���u�Wnѵ����!˟���L1*�6Z��ޫ����:j����,��BćT Y�����s�&Э���9��3�7{ }���8`�p�ek?/W:A�1�FR���_��h����!f�[�0NF�B$H��QMa�ޜHm��7���#b�BiR2�±��P�L����φܞ�-��Ҋ����.��������Y���è�b��1�YkA�h%�D�U���b��P�hM�-i�g\�V5hER(�̱?��LN�Y���7n3y�&��ǋ*ːR��)�o�J5������#Ui4�)$W_���;7y��'�?���u,��/���n���(��"�g\� !�3C�(|�b���+��e�J4*O@@kMX������)��gώp*et�&A��/Rv����o�6v���v]��V�T*�4e��*�]�����?@�#vPL'ט?�ϤxqS�x��"�����"��k���
%���E�؏���
�Hb�k�<^꺢��
Gۓ���$a���[ �m�s��8��^����D    IDAT<Z_w]!Jg��1������I}�3��k�iI��?}���lF�4�F#^y����%;�1�����Ni�(U�H�Խ�C��A�>�9t���홭��>l+�
�m���""���@{,�jT��8�\��
�������Ue,�BVd�!_Xt:�њ$(�����W8]4��ɧ\�q�~��������sV�*�"I!I x�<Ek���s,`�@zS��T4��Q��E���ZB�5N8n��f]�H\���S֝��[orvt��dēG)�����6J���R��OF�'��6`�@*��Q��3��4W�1�B�|��J$�ŷ'L_{������R�"t���xM�Ƥ�M�(~N���W�']���K?�ӂ�׈<�-W<9~��w�B-+~�!x~�׾���Fl	�}��혟����{�<�pk�%p֜�IE^0]�k|�1^�H��@�%K�6�iC@.AS�v����$'/}�i$�|�5LW1�"0?�!�G����S)|�gKλ�GWC4+�i�$�<C��yb��4���C���O��}��q`�Λ���/r�;�x�h]�Ĕ<�P�����!�K�Ҥ�iޓ�oݸś�hG�Ο�((��0������s,�N U�W�<V�(��u��Z`�� ����"����tV2��m�y�����{�E��P���@�e���C�%��:J�����)�M4A�ƣ=4�S�;� |�N#�������jG,� ��-t��#O7���"�na�`QA�!'�����á�G
C!��������!�<^V�&0��g%Z��&m@�ڮ%ђa����$����N4K
��:��ٯ�x�����&t�Q.�4������������K��tM���h��S��V��4C4�� x��<�*�2��d�!+B)��7ܼ�MS��C#(��:tq�)Q*�u��m@i�ܹ��B������l���>�tz���p�$k�҄� �7"�zvB' �,��_fpm�:�zE^���/qgC]2�`nVv��
=L1vM)���\�HR�/�~� ����D�
��5�C���!*:���!P��Ĵt�P�ܽ�.��8P��'�	��ĸj�m�a�,�ƒh���a��\V4֒H$�j��&JY5*Mi{���cm]2�P/*\0��HLcX-+�fs�=?��իL�SƓ]����NO�9;�Q��x�����T�:�#�4��ȕ �i;4���������Y�	m3#I<�4v#} ��|��� -4���Xw5V+�.���)������u���O����3l9 �vI\��G��Nȕg<�����',�(Ah[l�-"�2&�)u]ӵ�[���M�Bo*@/�Р$2�	�l�:�s�ܽ�����ë7��qr���O�ҭ�@ݵ��ϘUG$*0؟@����pB��H�f��ŊG�T'y�k�����>���Z�w2!�����[ "�(�KV�(	������LG|:�C��h-q��K9(XW�������;ܽ{�����8��d9M[a��q6��ak0�oCZ�$C��x�'hm�~�&�zU�5$YF9Ȑ:���HR��MI�d]W�=}Ơ0�)�y����"�
��� ������[����͝/��;S����w���xx����H���+���_z�����9Wv�N}#��6݇�X����+N� �������x�W�%��9v݀XcHC\�6�ᣳd@nO�!I��HilΒ��~V�l�H�q��K�r�����%$B[�A��h+��y���؁Y@�:3| ��D������^�xf��y92v��Z�V(�P�m�{#���j�=�l�g��_�d����p�U"��$��R	�KV՚R%Ԧ�s��()z�CL�4MC�&H�1m�m;������k&R����|v�cN��o���i���j:����|�i�AA�(����쌏�本�Z�zY��N(�<�۽�Y�5�}N\':�*IM�Ԋ�y>~ĸ,���T�+$�NH��qY�9Kk:oP�i> �c���bZ��DC���!�#��o�k�r���{�իW����ɭW���WHL���gsv�.�E��C� �`�m��w%5��lV��$�	����؅��Op��$*c<(cA�"��X�Nu�+���R	���:�{�[�	i�7�yJ�jY�V�et���v1a4r?�Ϡ$Jh���y�p8D�����^�㈸�᫪�Z�r�d�\�3�pxx���>��c;�?�Ç�����v6�Y�BX�p���#�e1���8��$�xHr]M,���
�bH����r�<g�`��tB��lPp��6��m��Wx}����L�|���4MC�bPF�����,�� ������H���p��".΃�4��Od�fy�b����g�Z�d�|<�zy� ����,%�4#(�-<�(�r�.�eA]� ��+�2��E�j}���{���O	:#_/ѹ�4(��!�Yb��9,��}�HM/�G�0.P5Y�F�#Q����[�mi�<�v'����tFq2��:��rȬȑR0ݟ�')ղE H˒`]�KC��[a#SW��]!��U �-2Dݴ�,�q6���p��`�%EQ�&9Y����G���*a�"�f�É�/K�m����_�w�[�rr�'�m���`��e�W��8�����ۈ���k轝��)��ܐӢn;��;vX�����Rj�v��Ϙ�S+���������C<�,(Hl/%ęwo��g��'�G(>�$Bh2������k��#(A4�JP2j��,[��qT�M�m�!E&D�i;�ÎB"c�҄��u���E�s�k��/�۔L����Y�J�&���وa$}"��Aq�8�\l�ó����D9IdW� *���tԝ'�:�Ka��n�B��9BI�T�)�qqq.��2����ږ\	�"�ZЬ�H�6B����ppm�������:���m�|>'Is�"g_g�r���S��<O�Y�>�h�RI�p+D�pـu�^��+��r�K|W�U+�<y�d4&�� �`�T4�.º�r���v�l�D���(�@�F��	L���dt�u���{�w��_�*n�9��G4�?��w������ii�X�~���;���A��	���-q6��m�/��[�9�6������^����������2�Q"���c\~�
��d��gC?��s*��ۥ�V�����<�zm}L��@����M����|��d��:���`Jp��U����7���YC]הeI���)�x`vzF���9l�<10MIM��c����ی.?c?��v���	�P�^G��x΍'sųc��Ox��Mʲ���Y�hgʻ�⛜�%v��k�zI�^Rd1	�|�`�Zm?�Jc�+:�N�������O���P!{�"�ˌ��[},I�D��4M)�u���'+
����z����W�`�&�e����*k;��I�ȋ7o�`~�OxrN��<{[���!W�=)�o֜��4u�4��;�����9�?����5���h+7���E��.�#:�
	��
L$t�$�Q��kki��;�y�z�f�ZB�OL�`P��X�bA%�$���^ܨx�->J�D����8��¼��!(t��e��:��^����Di��1�s��o�����g�`1�cl�1m$_%	j�0����W��dz�������;�o����[�@����:���t�`ox�k7_�Y��6�qz1\�OzW��r��Y�"�PK��dL�HZ�P��>?��l�@I��z��LIZ�bh����{���'B��W5i����h��Ŕ
���Q*��u�h���T'tkKY��U��Ԥ� D���C���� ��H6M�:�s/�H��i�'��(�3����и6Ʈ�˲��������c������&pi��f�B �En�N$�[��ZH���(MT"��-]�3�(Q�6й*��f%kgX5�f�C5_�����/h�%�U��
3	Hߑ�Y�\o�hR�鐻����kWIR�����3;>a6;AȄ�������[??�ѽ�y�яiϟ�3�XS���EJ͆��B 5^�]���/q���iۚ����Yq��+���;�`����?a�\P�KYT�,OLx���Q�H%"�xi�R"�scuG~p��o�a�r���r�?�	����W�ڷ�߾ŕ�ަ��UN<!	�L-&��C�^"�]�z��/?���lP��؇B�g���Jҵ_0����-k]k�^,���V�o��~kV#D��n�)�"z��D�Bl8˲dg�GQd�U����#/�����/D\/�K�1�y���?;;����>��sNOO��[y��{�� /־X���~M�'8�r��|4��B`��n,���d�V�p������w��1����̺����zMk�ۀm$�T+�g5E�Uuۂ1gY��۪g�Z��R(����՜���RZo�dD�)z!lC&;;XkYUK���������`4���ո�v�9l��9�(dd�e�n�Ÿ��d�lF$>f��$�x�c��s�A��\`����S�_���~��X��!cS��.�"�%p�8�W�F%	i9 )rd�P�'���u�#
���n�"t��l�^�����1����s���f��]8/���Zd}QY�P�\�#)G���l���9k)1MK�W����`��]@L��&v�>�g��$h�l��O?���?}��<�{�|��֛_Cc��
)2J��?�G䊰��������g�{lX��OA)ɺmHx�p�X2� 9Z6Ь���4A��i+B� ~���Y�|o|#R��	��>��u�P;G+%�mHw;;�D�L�lU!&|�R79A�Ԛ�YSe9���
��[K�Z�M���x=����vX�X��P(��`��ٌ�����Q#�
�2}��8��4 �l�v)Pb����r��d_�sq�\dOG$&.΂��Uc�=i���{#n\٥�,ճgԵa7��L �	"� ��]5%�E��,�w=�E�RJ��ƨa�`8���[y�j���?��Œ����k�{?�)��?d�:�Ie���D�%����F��X9�j:��{���8>>fP���/�"w޺E�eL�%q�r|��3�j����J�{9� �^���aݮh��U�a��A�K�g����r����YÇ�����Ox#mx���`o�w^���SOE����MDs�'�Q��E�����gm�/y��z6D��{6�r�H|c	ΐ���!��G�/��ݿ<J�q�Eg-"�8f,
�T4��vf�sق��8����{!DDv�$�8�%o���ɐǏ�8::b�\n	u����}D� /RlgX�V��Ӛ$�1��D�2�3&�߉����y���%qV�X}��;�p�5��w��LR�)�y���S	���WI���iJ(Lې�9�h⟈t;��TW�����ѥ�� r#��"���O��FU7����\.��PP-%M�!d�zݱԊ$Q�t@��U�0�ƴ��X��x�#	�k�.���Li�崪8%R)�ŀ6hN�����`XH��G2����Mٚ����}�v�P�$�4C����:��c�\ѭd�rr�i���x�p�aю�%���J阬����!ײ7��	������$�	�o�M�����3T�
�-i���j�D���zIR���	4M�
��yB�?k<z�ӵ�nI��,�8�{�������\��?����x�f]���dO��ѩ��ᇍ��Yx��b�'ѐ*��:���T��E��b#�����P�ؼG
�dw�:rwJ�4����i�E'�����B,�tuG��h���#�,i���G<yxJ����;��������Y/�`p�r:dqzF��	u��8��c���K�by|Dw��D�d���d<�:���+
�uMB:�!��舼�>���)o�|�-�v1����*�-y;�ܠ"���O�u�}�� �΍�\������sD��D�e׹n�H�T�Q���9��>E��5R�(ٕQ�`]�jY�M�2�L���e2�X�w�����������0$TmEil��]�����Ga��w���j�u<{v��~��ځA�@��4ֱ\��sf�3��h�S���1]�f)~2d�3��4�W9���h���O��Wػz;��ךE��n;�͇�A��#�]�RA�X�n�V���~�,������/+A�xhl�K�n��|�bց�ӭ�MՓ���:�yOJ��2f@!(�r�_�p��^*���]�HӴ�e ����|F�i�N�Y.����C��E���s�ޜ.�s�e� -b�\R����J$�$Jh�[Y���8��C� �!DH�uH�$��aB6(�yA�{�wnRO:,H����z9@MƜ��d�\�v5E=��ΐf�$�����i����~�Ρu�s9�6!��(u]#��:�"�(�s)mס���h�u�Ã+Y��$Mh���i"�kP`�����j���=����1+�Q�x�D�ܪ���ءKI�=2��i�����$���1�,'���Mן������*KQY�N�{�,��q3\W�m�Z�e�q�I�L<�y��YJ���}B�F�!���K:��H��ΐ(M*3�v@,�$�EM��v�Ld�U�D�E$G6uM�
���4uͰ(�4��ij��A��긳�p"8O�S�ֳ��Eҋ
��5�l�ɽ��-���_}�ӣ'��O���)&�7~������r�:3��!Y:"�+\t	�"v�P�|l^}ǟ$��TX��rT�ڎA���(�s�"4ޛ����z�H���f�:O9oi�
/]�u���&,e�Y�@'���,�4�Fh�����������c�@'Nq��C��?���/�����_�=?��?�N��ʷ���;�+?���|�ŧ��?s��٭�|���/�W�����Ͽ�w�>��r�����0�{�œ����4��l�yeO�j�rٷ;B��i�l}�`kB⹰�*�{�>:0���
�A���5pr�b>�bػ�O�3V�s�b�eֵe���i6�J�p�t0�Y�,j��E$��Z$gE�0;9a6;E)ō7x��W�Ӕ��G|���<y�������Rx�L�*	�G����}��b�I��%����p�3(����霣�#v�v0m��{�x��)��dY�i%���������;����|��cZNOOqy�h�Õw�r�={�������9�z�����w�̵_�E�8�-?G��1x�^�(ʵx�t.�³�ʵѦ�,?v슋B�t�/u�AQ��cR��{Z�Q�hd4P�"�],e���!EQ�e\�<�p�d0ܡ��mm��2;�HUA�b!����V�!���>�޽O�m,
��wFJ|6��Ey��G<��y�XgAl��m�v����v!K��$!O_��pQ�}���#�~0 �Mn��
m�����ت��> ym@&S�y���L�&%W�S�%�j�s�p"B�i��El)��a���#B�yI����ߗ*?�L�A�`X�Z.��$!O3���KJJ��"�H��:"I��iEG1�H2Mk�xL(��hT���bΎ��G���4���[�咦vtG5I��K��U�F�T����l�9���8K�a}����M�e�h�r
��H]���P-�;���i��U�ຘ	�:vL�Q�j����Fk��\�b�+6�R��뭌�E��U�|���AY��	�jIS�Y���1��w^}�,O�{}g�%*ф���脺��Ì�����y��Z�޾���0�P[�����0�~���\�J�e���(��B��񅈶��<����}��@W7LG�5���%j4`�j��1�6��6���gg���E(}(��k������1�a?nxY���SU�"%I�t��u`*Ǫ��p	�;;/9=�SgC�P�J�G9R�\ϟӵ-��I��p�lM�3���Kt���o2��O�0�y���ŷxt^���ɏ��ݻRa�>���z�����^�.�*x�l�c�xw�v����|��}$ynf��uG�i�m�R*-���    IDAT{ҔC�茗)Ks򜵐�`i���Ɍ����H%)�d:e�3aմT�p�W���;|��=�� k<E�3o#�!�2l��Tk궥5��'$I�3���Pu�3LG#R)PBR$��#��
.>32nZ[�x�R�4u�F�w������b�`4,�R��9�þ��f;��ѵ��s��oY�S�#���������C���~��+����0���7���� B@��;_�����+�?�!g'G(�(���t���:��R��#3����qo�����!�� �!�yV�5�<!M���6�2>�UU!G�A����t�BD{��[�V�C����q&_�5�݆P�YG����:�4���qHiHM��Q��?�e�y�oM{<�N�w�=R�H��dE�!˶e0	� ��H>8Fd#";�%Krlk )��.E�xo�y��ԙ����a�:U�E*�
�]Cש}�^��>��i�q^I���5�{��4V6�B�ի�=.�/Qd[XN�����
ʬL�Ʊ*���H..-c��=Ťµk����ԆMۂL�����gX2��ȺȪ�3�Ń�y������goo������L�k����͛�]'���	{��|�j��912���)2��M�"�
m�T�^�X{�z��YJ��#���n]SLj�ܹ�Q���C�2,�O�R��lLMUT�g��<�l��'��	�!t�vM���#��$K70T9N�m��S�X�x�'�tYG=�RG~�D�>�?��6)�gs�)���D��h�1�L�-�Ƣ:G.
����� ��&�<�L|�bݬ���QZ�o�H>��jB���[�|��PM�(
2�K��Tw���*
�e��0���e�����K�\�60�p�����u��KG���2�i<�4��E�1%j��Ww�o>�����_&?>���QE�.b�1�{��,��?�u�ny���8?�r���
�ir��nޤ�6!/BJd�R�IMJ�*�	�T�GzK�0�(�(Ц��Z�d
�. � �a�:�&mF�%J��
�����1ٯՂ!K�!�X'���G�"8lV0�T:m��B0;��d{S�NN�IQ2[bO�kyr�>���;��7Xv��ӊ{����>f������⣢;k�������2��:�#,l��x��us���O[V�Պ]=���{&h��C��8��u��6"�5��ľG������L(\\�D@�B;�0�D�DI�t���y��<�0�nN��W)DDjâYSL��c�Z�������w��Ff0t�L����9e�"�`R�T������MO�IA^�T�Qd4ޑ������m('j�yI��pѸIɉ���w=m�Aeh�6�v݌48�2)�!3%FGz�!���[t�]�AM�8|�m�pO�P�kd��h�X.�qP�(YQ_+�5�!��<�|mJ�k�TÂ�w�����C�O�1��c�w��c�$uq$�/	Z�.��uuQ|t����Hb�@x��S%�/��J#� WeM߰s��S�C0���2���=AE��D,q���k�dDt���;c�i�7Ivq�ϲlk��.�����w@
��~��1R���䥃����Lf��*c�^�)M�դN�q:��	�ƚH)Y+�M�N��q�@\8���2�������9�6���i����,]�z��oi�`'���K���ZI|$�o{K��������ՒfhXtK���/����R����WS�n����dǆg�眮׼��_ i���1���œ�,�)�$��G�u��t�"=�m��ﱽÕ��/>R�%ӲB��^3-Kt�aI��,����s�!&�fc{�gǄa�߬	�����4��G��Lx�n������-|���L���0,s^y�6/�	y��w�up�n��ɣ��L���/�
^R�F��˗S˼�8��e�ڢ�&�\f��t���Uhx������3��6-������Yb�@
���"���Р���v$�D�\d�G�v���YF%5�'HI�����c��w�H�
={��S�r-��2G�!��B^��ag��Pƈ�7�����ԯ�����*c-&�v��>���������;�Lp��T��!�/UI�O�٫���;NGcύi�R�d�9��D��YK�Z\�	x& ���*��X$6J���&%@�ٹ~���=V��o��!0��\���99>���)�����$��z�⫚�|���YY3�4Z���h[����r�&SvgS��|���v���0(S�xG0+k��������?�G������<;���-�����/s���,�c��(����H~S�|ÖQ��h����S5�X���V���F!"B�ӳ�m�~�pCOߵH]�Gf@Ha.1���IE�5|�����$�.u�#KM�X�S�O8���#��3��AF��������d'��b�~�c���X�B��u!��.�d�*��k��H��}�b��N�Ʉ2x�Ѷ�,�[Oy^�Y�c�!^x�xL1�����~����������r�����G�O�`������z�͇w��O���h��a(��'J��?�Y����ߤ�qQu#��I7�/��_�S��\3/�̶�TmRW�zI�!U(�Պe�o�#��7*�A��f;W!(�r�#�Akl�$�̒`t�)�F�݆�4]��bZS�u��}{!�����Lx%
��}9��+��c��'j���A�w��6rm��~yJh&�y�(*]�T�s8�EAYO�A���Yl��޻�ү��U���r�!@�<ē�=����ٔ/�k���������t���f��g�g�x��k�n2X�0h�3ݝ��(!�����ί�g�_�9��9�s�S3�kz!F�'zO�3vg3d�Q�i�l�<��_�:e^r2?�]���"��h&���7����Ӟw,?�ڭCz1`]I�_1?}Aa4EY�|q��Nx����b���"��h�q�Ft!A(ʪba-O�>bg�o�r�g�������گr��5vg��&���y�����?��gl?�n6�eAY�؂�d�b�BĐv��!�d�,������kJ�h$� ��|������;ܸu���Xm���C�Q�F�����&!����P��4�+��!%���g���{�'焇ϸ]L0yB���/�T��リ`��q��6g~����y�OcR��YXY�]B�J1��SM�TM��I���� � HI� E�"~gbJ�&ܺq��{&Qќ���K\�S��RC6_�؆
y=e��2�Xi�P� f2�ֵ�L
�r�p�ļ�������,J�.7�M�����wv�59������))ʚ���~���^Ń�	vZ��"Z�ě��Q�#U��Ĕ% H�K�[!cRz%q�(.Q"d�w/	���`LF"D�V�*�LsIa�1��"���@Ӭ��ۭY�N�����r6��$ �Appp���<H��[�[<���{���ut�&��1�Yh
-�F.!���Z�m����80z�S��ڞ;n&kp����5Ӣ�u���O�]/�J��{����ԇ��H�h1C��%�����Ï���z��\rͻ*�;��Ξp����Ϟ����ď9�	�tM{���Y��t�O�9.�$��)���W�W[��O�=B"l�G�9�Z$1hf4:�8>9c�܀Љ����� ����D<IUM�1��l��eB�g9����}鵥�{�<geҟ���,K6#/Fz�2:9x�����}�����=!�\�L�!x�L+ m�#����;���q���o�	/>�!b��(��TEŒ�A"��L+���ȫ��YQ�;Y������)��%;�)�+���&z�Q%�b��<?���R�;��Kv�g\[�v�9^ L�~ߠ�8?z���o�����y�z:���ݺ����(��1�x�b�t4T�����<ϩ��^�iہ����v��{wy�m��9������d�e���������s�<�=�i�5%3^�U����G?����[����S�\�f��oZBHT�0�DS�����{BjL^b��I�J���t}CU��������O�^��vc/H$>�R���[7K�~�1��|�w��y6���8?}D�9��%�^b�J�MtK���-R	|}du���m�Ӷ=�,YmVi1u�i��^�O��(]�{��ɠpk�;3�,C:΢ځ�������o��������������2���㕷������JK^��>�������IiOQn�+#���6�(ï���#�}H�t�Pɘ#+�臄1R���2���
���#�C�h�#���~��1Dr�Æ��?���>�^.�uF�Zqgg��޹Ba��B(b�1|z���̐-�����}3�a:�Ȝ�ŦG���Q���"�Y�s��6���C��9����������C�� ���5:g��_�ᳶ�Nk&2U�%�2�6I޲�n�)EF�y$�b�X��t�h}����_	�N}�	n\�U*'q��R���d�M)�fwZB�ċ�0���ݬ�%Ae��v�v3֋%��f�!�������ã�U���5��|�;����1��J�6�Y���(q�G�1�g\��
�B� �a a��CĈdW�n $&S�e�lR�Uo��	Mp�spp�B����|A�\"CR�w�',A�!S�Ar�����_�:��:d�������.{�N�T|������/s��_��w���)U������48���T�ٿ�x���'���
G�Z�ܥｴ�~�G/�X����a`%����/C�S1"�\0/���zg�~8ݾ�$O���,v=�G��[������8;9���%s�K�R���1�����MI��u ����yJ2t.-��2(Gl�9_���e��E� �8V ����9u]��&�+���B@�nX1lZ��5���ۯӜ�"�ݠ�|��ѶL���g����x�UZ"��B18O^(�� �v<~����g��w�w��	��	�����2�2Ec��-+
"��o���?f��KӵU���޿������!F�(v��)�Cg7@�7tbY�$�e��'���r��to�|R���Y�����5O��ǜ�W�ˆ�j}DK�:����"��9c��]�(��a��VoUېN>Rʔ'>���J��B�d)l� [�i�%��f;|��_`����Ɋ	��$��*�*�+��b���vx��@
�'��>�����Y.N(&Ez�L�����J߶;{����g��7�y���a�\���p�^S��?�2�����Y��.� �eFU�ɲ����'_�ѷHF������_�#^����)�nI�7L���H19�蕯rx�:s���s��?�s�^r1$�ڸ)Vr����I�� Qe�цH5a����;�P���Ǉ�B&��PVȼ�q�� ��dJ�bD{h��wh/�rMT���j����6kr�F�M�.Z������%�~ ���dy�e�@I���8���y񂈤�sJ#	~ G�>F��9�����4/8;=c���q�G}B�zJ�|��_�߿�9a�,Mߠ�H=�q"�ΦЍx+F��*JdRI_����ޏ��N�/Lb!��H��Ȗ�w1���C+�S%؝$k��'M�3O	�<�j�ݚ��Y=��y�c0%��8�vD�3e�{HQ&��jq��y�q���>rvv�u~��1-�C���X�_w�#�d�Sc_UȔ�1V�"-x�X���6!��	��d�~��cĐb�sm�u��Đp�1#��J��C����c^��_b��|��;v��3:JѪ��W�絷>��Y�������BŐ���g���zI=�㶴�f�+���O�Ŷ����{ReH]�޷	���	Wl�ɕ0l[G���>G�n"����|�y��&��8_�B��/��&�|�-b�|��s��9���@�'�|5��w����k�m�r���r�����"Q�V+�L�4���n��
- A�dD�H�`�\>0��b����pyA����9�����b����IB��Fbc���s�O�r�?�^Bۑ��#yl|˴�0�TY��0�+r��í6��s>?�����|G6�$����`WKT�RgY�]��zT�>)"�=�0��;iY�=GJ�ُ������yA9�Q�S��������$+rLU`����x���H�AW�*�m�}�3�z��r��4��{z�������lzס��[+�|N��赛�z�z0C�i�����d��:ym)R �8����DF@��'d��w��{��i�Ⱌ"�B��d2b��������=�uv�ݴ��'�~�b�6+l��TEH����8�������a3�����[��󓧘B��y=a����5*o�ۆ��ǜ.>g���<e��9�9��f���S���q�Un�N��	O���g���
6��:���{wy���k���߽Ϗ����	Z%?���M���v����xk����jֶi*�BC�yE���W�0�>�
d�)	��;O��>��%?~�!��1��.'�AѮ��eF`c ���FIC���;K��8M%���e�v��=�v�z[v�!�2֍m��n9�m7XAj�d����w�.��� !6xĦaz�h]�4>P��K�a�S�ܱ��yDs�L'X$�$�Ks��j�>�vf�W*.�_�21:��0�h)e�R��BUS�uPt�"�H1ý����=��P�SZ'�J���}�bR3��FU����(��,���_��_�9w�ܡ?�������~�&�sb�m]%��0�.ӆ@ �  ����C��f��x
,Y�]r���0ptx���h�pI 0Z�KM^z6��(�{�U>��o2�ȣ�}��������fj`>�������k����x�k�?|L��Q���BIu���ӯ���i�)����9� .�$��������4����z��@���ߎ��G��h\,�&=�V�-M4Ƹ���� �����[7X,<~x�G��`��(
�z��(���Jz��On�i]��?�U��x��>�͂�C���v1_quч ���{kS�Q�ԇ�EK��V=��1�9b�d2��Mƺo�H��*/�OszL�)���YRhA9)C�Q�b��?����{�<c�^"�����д���Ү�xg�Z��g����2�&(�&���N`�� q���>8ʲd6ݡ�Z:�R���G�(�Δ�u�|�Lj<ѝ�E���Δ�`�[�����i�������+2)D���ap�#W�A�
%�7�F�]���U���4��/�I���𨻋r:�C=ۀ�@�c�IY�,-.�%�`�A����4L���}��%�9�!6���F*��)$e��	���OO؜s�\0�n��ۆiY�E��$V�a;1���C����x��o���z��)m�0����]v����g{j��@W�e���MA�˔ 5��f����|��|��}��P��ǜ}�G|���5o��z� ����1O��m^y��W��}�7�k�x��$!"b@Ȉb��M���,�. 1=F1$R��0�!����1�:���h��]��(1¤��T��@�R�F��#��eC,!�YZc��rS�S�sl��p��܀k�8S�<74]:���dfP&�]-S�A���\f�iA�uئM��i�Ԛ��QH'�r�1�͆���
^�,5�&�4f -��1%���~�ڂBd��eL�2��P�C�����2�}��� A������H����>�Mj�4�3���'�j�9�YF�肣���v�6�iͺmȲij=�l6���#����x���y��1���{���ہ�����<l��i2���6�)�S#3
!c���d��Δ<���	�ł�|���	{{{�Y��SǺ�Y7��%�i��p֝r�k��AnPeΤ2����������4LKA�:���9�7��'��)s���>~.KK�߸��,
���\^����-G�5޸�]܏�ﺲL)AQ�����B�qc��ڂ�6��g�5��^b��+=v!�n���͛87��~���I�)�j��&������OS!X�V<}x���d�7�|b<^�~BL�<uы�����R�2F���6���3    IDAT�#���Cg�F� ��CM3\�Xl��(��5�Rc̟<�9���y��=6�������X����f��0��Ɇ�E=���Ɍ�����BLo1�e��F�(��hi(��]�X��s�IL�~�IB�r��;>���VƄ��*��I�+gZQLk^��3�a��sN1>rk��:/�C �K�<��]�퀨���B:�`[BY����Ct6H(&��f�yp�!�!���+�u�p)P$���������@�c��m��gd�_�񽻼��c����Q_?"�Mq�a��X>z�G�->�ַ��9ZD���kT���A�*%�� c"L
���Qz�S��'6��̐*�7��2?>ey�1�� �nY��lo�<�u��Kt����L1E���ܾNQK�ر��{g�i�>g�|�kŌ��U�����}L3�p�×9q�W�T~�T��1��Z�e�GP9���\8�{����nI�5cFI���B��
0�g�2'�K����ʓ�ӶM�$�r�&���#>F�LH�`��`��(\J�
)�Ʊ��s8g��"7��~[�̔�.׃��:�U~���&��}rAL&6�%�A�(�w�L#Є~`�l����r��b�@�!&d����=1K 1&s\�������V��N���~m| �H!�*R0���,Ӭ��n���(�(�}ץx�iμ똾2cg��w������_�9M���2�v�����M��w��,V�m�R�2�)�,�q#[��VWpebB�BGQ�e�}�6�@UN��rrrB��5�xⷴ��n`�4Bk����'h�A�t�=���S�32�9YoX(�ΐ�%*��Pm��y�`~~�6#���jtk���'�[�����r�'��'���B D�O�2�>pl�0۹���EW6�Gy�@�ud�F��!=��g��\�8�gY��q/Z�α��������z�6J�����`�u<}������}b��x��M�Ҵ=�t���>��v)%��pA��ap�o��R�6@/;��O��d�ߎC�F�&4�$�U���C���\lo�e��8��4/���~�s�G}$/+��#ߛ���U��Xω��7k�~`�]"����6H'�^b���4�ki�h��=>J<2�������Za�	ߵ���|0�pAx��N4kix,U*�
ϑ�aS���y���#B#�k�f2�8t!�B ��@ָl�xn-1Eq�Ǐ�q�QU(�ru����6��@�%ꝓ�b��UF1�C��{�kYFK?U{�}:�̠���'�������c�h]f4��z��l��t����@��k:��Z08�Dlm0���)l�%�L4�(p�a�r۱~t��8���%+d0t����8���yF^�Bc��w��c2�����k���-Η'�K���!�����\U���[��	��y&#���u����4�9������@@(A�;FE�On-eb�K���c�9(�Cn 7q����a��)��Uo��f�jT֑�7���.2�H���SBH,ta@���S�9JA6n�Z�R�.��LJ�"O��n��20&c��ɕU�G��#$����:|!p�"�@��JR��B���>_q�h|"��QZ3��5�w�9��<MfpDv���%�~Mɔ�;L���Ð��(�`dD+��)PIF���d���8nk�+F+\������4��6]lh��t�k�>�ϧ�o�^��7!/����ES��凞�v'�]��೻H�y�wY���Y�.05)<;��vD���u^$ؗ<�+PYI����CP�6px���}����y^�ٖh�dQ�2Td��I����!��JCA�\�֣ª'���	յw9�6,�d�3��v��֫Մ��:m�����d&CF6�ֆ+�?�
�R�~)���S1(|�XzO�� �$���V���e�2�����`AI����1t=.�ZbmG��1L&q*R���>S�0йm4.X2	RE���a����$�sαi��6�2o�Q`�K��Yr�)��v��ιq��Ɍ�dB?LgYQ�Y��l�j~�b~N����!�j��B���H�L���r״4C�D�uF�NE��i\&01q�e�# �7�Q%�C��s�@�sG�?%�}��������s~r�t���Mn�.1������]�:Yд�x���J����F�r�֢tgΟS�Ȕ"�`�5�`���o���RH��c��wc���{Lo�s!5�t�jgFV��� ۖ���
��+|{��K����8��%��ͳ�3���r��>Eb�a�)$A�4n	���%�2�K��Q޺Mp����Q�LQ"�m6���{�|艡��[�w��P_?�>����1��:<����C�]m8�ڀ�փ�0��BM��Ve���E�HB]`�@4�Tl\K]�{�X,�s�Қ�[�מ�/�^�'3VN���<�Q�+&N�G����d�1e�λ�V����u���-��2ٙr~���{��j�����\�k-%��T q�y%>~"Z$�e�2�,�A&UL��(5�[$�AF�V�ٽ��
���5&�(.���s�<������9�yՊ ��Z,�N^�Zڈ�yN���\�����>�T�W��?�7�'�2JfBQ1��.&/֖�v�F�d�s�`�Z�>��ӱ�8�I��R�kݹ��aB��Cj(�JH���E�ϳT�������2���|u�G�OYv;���b�Xr���b��Ԥ�,�"~����}�s,s>���9~�9Z�dF�t�^�Nc�zCn��EfG�va�{��������l��s��&�7��n<�z #ŗ-��c�ko�F���Z��'�ke�,��Q��������?��_�&����7�y��<?Eَ�{*Uq��� �g���3l�%�MHσ�����?��ie��cn���0w~�RJ����۹չ�>�/^��w~A��1��r��D����R%/���8���)B�2�t:�Mi# C
�j���H��z��V���4]�67Ҋ,�*�m��w�\B$H�*ac+!:K��S2��)sd[�T���K�c�wb�H@���0$O��W�x#1;·Hy�Unߺō N�L�g��?�Y����}3��,S�}p��o;��5�b��c��ꌙTt�\7�uK���l��+�߼��)������͔"�@��>cdR�R�V��d�w�tg]��>?�'��,(���-T��������D���l���rC!�Nf9�h�>q���m��������j
ȯ���7��������Đr£�2��Y���e$��V����)�[��R��֊>X��7+�}�!/���"| ��Q����x��� �L�F�|��k�L-�(��C�H�w̐|���<}���^c9?gRܼy��zɭ�7�d���ٯ��\��W���������y>���a��6���an����v"Ju�lw��������w�ѿ��'�(w��BI��x�R�3��}ZąN�-.^���#S)�B-������w�L>�����ľG������TR 5R��!Dr�GL3�ͼކ9��U�^�%�K}ő-��\mk�dϺu�t��_�d������qǲsν�3���F����mQRSg5vpa����2ٍ��؛��%��r��^��F��O�X�������!D�����s����NM�I�!�"S�ϟ��{����9�����'4��ǧ���Ą�
e&�h˚pp�p>�9=���\z����b��v�!�+��-�ږ�K��l��e�3�<�	5i$�L�w����@����-U��s_~��y�X�4-J%T�r-�v�Bv3���������x헿N�7��sjc������9���=����I�ٔ�/]?��ű�Ӿv� ]� ȗ��/�̾8/7�i�_�]_�T\����yڴMײ�;O��֊�s���򒮳)Q5��d{`���M�Mn-s� R�hR֊sE�t:��:��iZt^Hڡ�X\%4�z��j}�Փ����5F�)j|.��㽸̙��ߗ���*�������E����u��L
B��|���!QDB���qH�M? �B!�Ҡ�&xI�gk)2��5�`i↮W����`q�K)��N���:Kc����J�H���!��*U����(�
�d�&�UUSO�(�	*S�l?�ڭ�O�A�:E%v� ���K����d��})+��$����(�u�%�unX=y�p���'l�|^������$2|0�q�$�x�,,ro�+�]��Yl�!�JV�9Y.Pr (��O����k-m������?�M���d���%u]3�ԳG�$�)rڶ��(6��:|�_��or����_�~�!�o����.��9�bF^LYt��|�'�g��	����O������i��ʗ�A����dX��f|�������؇�q4�2�����M��?[)�N���')��5F��v�̍J"rC��	�[oQ^���k�4FR*A��"zv~����,Yԉ�68\tTe1Z�Ҹ���b{Z������m�,��%��&�ר$�k����z�:f_�B��M����c�0��BH
�/
����y�_6�[v���o�q���q.J6���'�u�������	�*Z*�wcO����Ag�:r�s�(v�	�4dY���&���p=|������E��g�x��1S7��@-t~��p�#��Ͽ�_�%��kt�d mǦo�MK���0�FѴ-&�b޼�ɳQ�h�����04Ӕ�=M�p���f�lFx|���Ӈ(I��ABg�G��LX�M�~���?k���?r��ց���"��d4�c��~��w~������ѓ%�rL\�����'��_�U��j���gT�s�QU�ґq�c�a�/�ɤ�%�M�ӗN�UU�`�<!������Id:�R��ݶ��\eY����\���#R+���inݸ�믾F�4,�K<۶�(��-�z���9���J�6�52E$�b���\`�H��xA�]ZA\0�K"}Ak�Hz�ȴ@IM�K��r��ЊvqF~������9��۔u���؛�H��g~��|{Dd�VY�U���R����DR���� ��m�ط�����a`�پ��a,�D-�Dm��ޫ�k_�r������դ }@�2�2#3#�w��>�ؾ���������f*ӷ���Y\��'ۺƶ�m�����	y����	��3����$�)MUMs���cuG�.Dq��a#��2�PqB�dE�hg�>t���r�pL��,"J�ާ��T���3�s3������E��:(X��,U�dH�IL��/��W׊�5I�[��%���?su|�ۿ��s�i�ȭ���4�z�EŢj�s�R����9��{�qrp�m-Y�й�4SD����m���wd:�5������?�K3.�E!PBFj͔-������Ǉ��3�+_"�Z6�"mz������=����N�G�e�|��`s�2ɻ����'du� �?���������"�F�Ve�bo��<y��?y��*�lЙ�]��w�:�.djGJ����bm02�xܲBw��/����B� JE��ȥf3�qY������OnS{����V8)轡�-i���5!������M_�rXе��$�^8'��l�p i���	f]A�����������^�e�g�9�u g|�_����W���FGpt�C�~�'���f�P�g���e�IU�9�/���G�0w���P�n���j)���0^ctD�:��8�!U.�6=��8���������Gwyx�4�IT5��[������ЩY��J�<~F]�am�P��uI)���ҀN2�����TΒ�6�k�<]������R�Qh|JIPxK@���i898���a���ZGHI��,�A�<�����r���?��Q\��@$gG�f
�i��Nf��);�-n�����\h��u�a�bm]\waf�U������������U!�!4+���$/\]FgY���q�[�$��kt�q������<mFq��������Is�� &��.fz�֭�oǣ���QJ���SI��C�cw�ܡ�*���;�ƽ
���{�+S!�@إ|��
���xͳ�����!�`.ZR<Q��p�R���I҈��'�D�}~��oB�e�4%�.�k��P_��=ASk]O���1��إ�����\`M�="��uG!5�$���4�:�j�X�#"�W����RR�'GE��2�8J��`H��b0&JB4�P���1�����Ɏ��ef��I��t�%;[\x�gn��Ӌ��B,���bI)���$}W3�9�����c���V)f�&��(�IV8�r��F� 9�JH:�S�-��f�(9:xN9]�����9��"UT�)�p��S��5<��{<�s��K�|H��������&��ᵝ����-ʶ��h�O~0�����l��Ï�t���;��y>?�:;���������jF}p�~0 ��=�5<�%9��h+�֚�FFU�x�M�2t ��^I���D��j�=oBjb0��n���5����C�/�-��0"���I:�c5F��<eQ7(-ѱ��z���!�"���dY���MU3����l)�{�������D`j�i���۱��.���,�/�X\��C���re�)V��b���֢�!����Cڮ�Z���w��?]�'	2N�:��8Y�$ŀ������b�l���Br��=��Ha��Bi�TEc{z�q�b1�D��j<=|����K���|�uT�QWU��ZKo��^��(B �b2��`N��Kv�!�	}F��q�HSM��e�9���gDZ��K���CQ��Ӵ4�'+r[� %�ix�ZD�b��l8b�d�����7�dQ�"�3"�Q�Ϩ���х^Oˀ����I9g{0����O�&ǴiƖ���n�AJr>ST"Xa�%A�������&�}��������?���>��r�B���w\��cZ�?.���SEx�XT����7ߠ�~���B�D���麞�d£G��z�
{�;D:aP���Ή�E�P�w/2s�r��]���)5JH���YY!�g<�TD���s�J1��Bb/M��LP��$���J��E��K1�E��ۖ�jЛ����7ٺq�����>c1��E$��{�&��:"Orfu8ꮽ�g���,�ԧ��o�������TmMUUP�,f��!��$��ic�h����#���jM۵!)HzV�R(���t�4!]�G��8�Rc1Xa�	H��;�tZҹ�.H�׎͗�z��B�r�^l���5f����c�|�;t�a@7Ӝ���)Fjy ilX���Itt�1��8
~u��v���YT3�yAd����Cu�V��6�/�:�Ђ8Rt}Eߴ�Ռ��FG�,��.8Zkܒ��Iw��߿�����s�i��,�������]f�=������1y������mIi6��r��qJ#�Ɍ�ȸ�r���8�ġH���!A-����A'��IQ��X"�QB�}X��y�r&���/�:��j�F��qV�$C�ӜQ^໎�y��������s�R顣(t����A�h4��w���ի<z�w�2�L�s����dc����a��뗃�.�͋���y��"����/\J��Љ�|8�P����{<9:����8�˯��JՒƛ����pV�`o<b���{!II�e̒'�9�,K�℈�Ak���8�'�%�wt�	�W�s���Ř�HK\�S��E�Ԋ�`#�b�C�)��3�3�<	��3T�s��sԶ�k�gg�<����+��(I���._���3�v���`<j� -�!D
��-+��3"W��g9q�Ӷ-'��̧ST�)�o$��9�Ɍ��^��5�29~�u}ٱ��S�̦h��(�!
<���"���	Yˎp5�Y��fG�"�]��/���
*��C��!K_�����V^$�����W��n~P���R��
�)g@8`    IDAT��!�g���m���23~������ӎh9
H����W���b��֊s�����<���cL�A6���i�<����h��dB����^,��VϽ��Kr�U�BJV�����Ձ�A���G�-�,缮i+���?��;dv�S?�7~��]���O��������^g�4$I�0G��s�*K�tD�br~���>�I���U
g�=i7?���+�����m���C�Ƣ������wo��w	g%Y�#��F8v�I��X�ϵ�D �@y�QB��р(�ıy�q��bd$�M�-�LI⍐fT����O��O)|ƪk��&�Vϊ&B�����{ּ4��a`r}LOĹ�q�������@�G�FG<��T`�fqf��cL�!�$��m�#�3���1�(�,fT�)բ��e�%R�'y�"���cA�O#�1y� ]�%�z�"��ֆ�Ju���W^�8;;c8�dw��A�9F"���%�����+������p�����,]S��5�Pf2C��/�Nx���������-=�����uS3�EJb�m��ՁLh���Tdd���1ny�Ǵ���,��P�nSu�4%�Qňv�`� ������X(v7��(
��¬�7dJ�/=��,[V��k׮���G?��K��Aü��l@~��KҞ�iB���v-+zis^���~��/wT/sL�x]\�>�&T��Y��_��M�����pew�G����'��!Y�C,��윃ɔ�(�q�*ۉ��s���$��Fx�]GgA����Zp=�� Kc�y�1i1���i��/�S�UG��1��>��}���.�i��&Kr"�d�@d
��C[��q�#�C�LאHM�Z�v��p��í���È�y(�c��x}��I�8Q�W
!B����-lo����i5���'�늫W�p��WZס��wX�5�Rxkq��)��hu��5��[t�5�Â�VhȲ.���$�.�g�L(҄B�X��c#!~Ev�箏��������Ϯ�/~Ϫ��鋦��[��\ �	�����v��c�!�\�;i��̦ܿ{��ȉ���i����)�-�G'$I������$���Uų�O8=>!Z���qLoJED*�/Fˤ��l�`0 �(�*WM�p?��Y~�ug�P����_`ݯ�{�[��@{lS��5qs��`�%��tP0`A��w������$W6�5:����Xe�M�(���x��4������"e���"�L�8�MϐQJ+s�s9͹��Q����C�L��&�	��:�a*Vi�R@6��$Kb��Ʀ7�(��A�(+P(�,#m TLEha�C������F��o������h���p�ӵШe��c��'׭6�ē�HC.m�ಁ��$�1�`m���������_�"2D��|Ge�ӊ<+XT%Ÿ`Q��Zp>9FyP��l��x�p��t�SNϘM�0�g�L�'g�E���s����ɂ��Ì���y���^�w`'5j�����G��"[��{y�ݯ2m2����f�T<{��˗�y��kLΦ���3��DOK�>B��Ӗ�?�O�݄��~̞P��;��d��;�~�������#������J�~�P�г&Ġv��A�LN��U���&2�@�hk
<i*8�:j#����餅��8�!�CHŢkH�?�>9�ѤDF)���53$~0di^{�u�����T�4�(��*�(��:��9�ٌk׮�X,88|��
-�Rfx�[���m�ش��{A�#��)��Y�Hc��3=EQ�4MH��EA]פIN�5(��25� 0���إd�X���|�y�����fƲ�[BߑҜ>{���1�x�?��;���=�~��rN����9"�y��e��qzD�D�M�gX�Q��Ӳ'�2G�iq�g��S�1s��KC}2��=٠�v5�������G�v��kWI�!'���|Uc5A��A4*ȣ����j1�;���4���㽧�mբ�.�}��m�|rJu|N���Q�c����O���tޒ'���`csLg����渦�3���G<��Sn~�U����x��_�AD1Z��`�B]:!S�t��G1��pI��N4��Et�(Np��Mc��O�DEA�v蚆>����_��CH�Z���1�&��Z�}��n�%r1�9���`�GE	�W����QBg+��(�C⥫QV��m�A[�0�}D�z��`Lp�Cy��AJPĔ�!pض!��~rvww�2x�;<G�D4]�B!�BA�ft]�J���ْ/#��ix߇��8�֙J�~>����`kg�ݽ=�OO)����i�'���*�0֓�;"�KU�s�#�[�8G�Fsu�/����nB�Y�R�X�o{�KrWm��a[�>{����_�F5�Эe�5},)���j������Ӈ��ߥQ 6�8��YQ�x�2����S���3-��0;|�sg�v6i�������z�5��Ǜ�(��:b��0�ZDA�8H#F:"�"!8t	��E
�����&^
ـ,I1⌤w�k�I�^Af1�i�\`4�	�����g$��C�A\U�A��r�}��_�އ8YeY���-=j�Q`�)�5t�p�e�4&
�D�g�:��􎪪hzK�&������qO���U[����&��6(?y���4m�m!1WǗ��y����=��bF���]{��K�Yɐ�K����[4�A��+d�\g��I4�@]�IҜ���bv	����go�{��g�2i{���m����0�r�EE<���o"�7�տ���_�)��=���}�{ޠ���o}k(�Y�����Zǰȑ�cR�)tF��kz�	Lw��ޡ���$g�ګ�"c0*���������	����ɽ��<I�����b�u]ǣG�ְ���y 8"ְ��`5�_,!�e����W��r}ȯf�EQ��z�]��4M��

�p8�,�˟-0�ǹ`��PUޫ@Ҳ���+�~6����wvȠ��\�s�Jp�.��
_��*�o�?��Y�H�(�(1��xƢm�*&I�S���|��K���!�Y��UOU�0�D�!��T���Nx��}T����]E��DH26�G'*ڠ\,� Gu��JQU��/�&��vđd#�puE?,���)ܴ����C0J�;6�!��qI���4	{j� ���%r�T%<��!��~��-��6���d2��� �b����7,>�˕������a�%BA�	��ȦGws��4��dE�Z2���B�l} ��pK��������_J�݅P6�0�'�
���Y?���`�������c�c�AX�}�$���Cv��خ�����J��c�$C�u0;�
�(<�4+t�P��f孻���nܹ@�K�du��foo��bA9_���{��M&,�����	�ąl�����9O�wƗ/�R���z¡/B��2���f�>�s���?�{cҔyճ�w�^'<�gă�"J�yN���ޑw���x��{���R�l�x���������u�<��	?�������U��t��tv���%����Y����QR�୯�"��q�����矑N�l+ʹ7Hy�r6Һ�ES�ƚH*6�)�	���;���1q�Ru8OJD��^���T�e@� D.�?��g��*d�@�&xc�
��tN`��i�����x����!�K	�AY����{ϏPQ����U]S�5Zk666pU�oڪ
3ʺ&I2\�s��]N���`@�Y�?�����(�q�Ķ-�|�`���لj^�s�2�c��G�yp�t4୯����.��v^��5�E�x���$gZ����N���<J����>׾�_P-J
#�]��&�g���\��WQ������������>v��
*�0Xu��6���XcKI�RbZ��;����t�J0"��q��w �l���<b��>ͼ$�
��ڷqՔ�yͣ�Sd��P!��kZ:�/;����cf� ���>�Zn����`:�2��և��,˖d����{�<�C�X,.hw�uW�eYx�����j��u�I��^ҵ�:0e���配y�!�b]DHB��`k�o��o��7 �A�b�'��c����`�bs��miNQ��AZ ��E�r���"���{$=�,"Q)���	B#}B����e��ۢ���z��/q��/C1��Rbi�Y'�	>R�2>��tm��=m[3��� ��eE��8���
�o�gz):X����
��t'���12M�3����>m]���9V9��<�)�0�*�il!u�iE7k��%��)CZOId�QI��з�`.�
�F	:�1��$�	`�k_@����ř���K������r�z���� ��y�j�V8'�횕��A��9�"m�29ӡ�aT�L�����[ ��$���{���Y(��EmX�t�ǩ�I��a�w�E�h�7�7K٪8_�+��{�N�{����4����ρ@�K�)4��PK��i�
���vĊ`��`��ř��0Z(�P6@�\���w�7tI��u�2�+;���\���&U9�_��W���_A:A[�|z�3�ݧ�W\��d^�o�3�!���X���[||�.����}���#b�(�����2�R��!V	��=���L��Ԧ�"a��k�_{���6�u'��B:~�V��6LS:� gP�bzFy�iʎ�u�8�lk��ش�����2�_�刋�*/kHY�}���ª�UG��7xQQ�!=��s~��D��)*>���1j8���>ۛ��}�+��c�����q~x�Y�q��	�O?���sd�#���nQ�^]7��.�s�D7T�)�>���
���<��k&���|�A0���ާqgyz��(K9��=66�RE�hGhz��cE���������׮���_ď���j�"�˘N̑��v��M�ʑgr�u-�qt>b,b&ˍ�8:��^;�'����{�9q���ۣ\�Ֆ���L���t]�O�{�J}���ì����\�0�9x���#�.xr|B���j�ozi�����8^�蛦akk�W^y��^y5��ʒ{������������(��׾FE�eIYιu��ł�ׯ�ꫯE	>��������_�����LǼ��;\�|���S�<y����ឧ���k(q���e�(_PN�ˤ�U'p��>���L�g�I�ޥ=�gO9��6f��̬G��D{Hbf�s�5ԵD��D�� %���-ie�PF�4�aV���R���'h� u�\x.�W����#z�	F^+Rb״a^�Ĩ(�7�ଈ�k*��B)��=m�PNgt]�d6�3��,�?y������B`���w6���7�w��'��x-I�<͠3t��d9��>���ͯ�ŵ�{���Q��
M���ofO�a���6&��G���?���6�<gR7TQ�V
�͉∲�8�%�J)d���o���qň���;�/fϯ�����!֭�J!��D� ����/�X�ڱru)�R���� '�*�nc�RYk�[��	��JGԆ��QJ���8����:����VgHBs)U��Yv���0�@�]�?V����ڶ����R��s"-��!~�R�����2�2b5�>ح��a�Dg�/^�U �*=j}#/I�^���_z�����?<��	�р�\����Ư�
U�o��f�SNΘb����+=�͹��;�C��̪#,�Υ=�-%�ł�tZ0�#u�Q\x{
��і��	?��Cڪ%W_!��f{X`�	�-ޓ�r�.�p��>�<�s����+ڇ�I�Q2"�k��x� ۉ�-E�!�\/��-	O�
�/dNn�)g	M-;��+TRd1�����o�{�7��]�Wo��ƈ���������ѝ;TbH�3ؠ�O�OO0�=�W�T8k�G���}���`�gx%�z��YΑ3��ڑ\�c�������Zs��]<��ٌ��Cv�v�ڲX��N�t>��l5ἱ���_B߸�1[����~�#n|��l��T'�]O$<Z+�����?�	�G�����L�= Q"T�^^�J$R��p��-��f$S���7�mQJ�=J�*�ғ����.��Y�l{���=��a<�1)Q��d���x��ã�܍�xz�q��]��+�����pȍ7�N�y��)��7n\�޽;(%��uM����\�z��w�2�M�y�&����u�w~��!hۖo}�tM��˗y�Ɨ�u�V��o*�j�[o�ŗ��6M�0\g�2�g? MS���o�����W�\ᣏ>���0H��Z���n�ݛ>������\���D���>���)�iD�E(E'���8�'!A)��5dw� ��6acS1�K�ְ�MkPR���ǒ;&������.�����Dv�yD9_�� Or�,�>G[ͱq�� T�w��[���Ԏ�x��8�c\��=Y6�ҕWp���g�ќE�C���*�^y�eTƠ��*l�2ր	I���ls��e�._#�7���#f�D#��:��4�aB�s�5��}Zbz����3t��l�\�s�W���f��ϵ�}��xm��E-�����j	[�BE!�j�/�2���
�_�?C�_�f��	�� �5Z$ĊH�T�x�v�b�8ia�߄,
�%B*LGŀ����]F�C���^�PYQ�> �K
g{��K>�'�
#�������@�̝����AdKc���B��^��\k)˒tsL����y�B��/!|)�R"](:�R�%|x�׀�� ���_�.��X>��;����x4�J\��:�GC�����/)�D�7!$&%����SlP����d³�3���PZ��c-7�^�*99>�VJ,���Q�Z+t��kI����4O��w����d*����(fsc��
�t���ټ����6����l��~���)M�gZ�2&�z���@_JP��xo���K���8���p_k�C9�S��AKɈS��`�(�t}G״4MC���8��-#d6b�����M�׿DO�R�!�^(ꦦ�{��M6߸���M�'�9t�	·$QB=��u-�C��(���ΣED�3"���X�S�K7��o���}�g���%������%{;�H*�T��c�'�Ov4��k2� �Έ݌������ ��|��ڗ趷��	���O�r�o����-=��)�=ZxD�p�R��-�Y�$�m۱���[D���f+�����Lx.E"@�|�[�?{@�#�yI����I$ׇ�s���g��Mn�ʄU��Z#q�Ya�������3�F��_}���� I����ߧ,Kn޼���v���o��ohۖ�}�{�q�����������Z���ש뚿�˿�������lmmS�8��?�	]����~�$ɰև�~�PXmf~I<��`���������R��O����3�'O�7���
�D;h��6���"�Q:V�Y��0#��nBN8:FE)�aQwX�t<�
���T��}���"�qDt��O�iN#�y	�Q�����R@g0�29��u=��o-I�)�E�:o+lﰋ������@6%��Cb!P"�"خg���y	*e��ʠ��%!��1��'癏�$�$M�bL~<Ab�`k��x��l����G�$�&n��OS�������nL2'o����~�*����#�����7���&�����n2���8��?��O����������!B�����Y6���/Pϋ��*�8�o	YDw��E2��[�W���RQ��5.�5�#�|�R.4US�M��1B(�5�}�$��fQִ��	g�A/�(��|��P�%�jm�s�#�U+4a�����L��(XK��4Ib�%I�p.D,��^�����/sb9�]�bi�*�������C�CH�"d[{�r�l%
ml���%G�O8:;g�����aQW�e��
�(�t;,�����c�����svvƢ�3�q8��g8�0F`��B���=����B���I�$A��$M3�����hw���xw�l�з��������������'��1�Y� �Rt�@VxT<��nkA�*Q�2Q�Y����Þ��:>8o	@� �#�%Q�yU3�d���Tc�.�s�שN��D���z�t:a�ꕀ�8W�0y    IDAT�R��xr-Ȋa5��h8<j���ls�f���çtUKLJ���H�b�VE�v��ބ|j/�2b����2����_�
��������e��"�2E�dzF[-8p��waN�,*QX-2b#�� ղx~����8��#�������U:��h��ʲ����E�@���H2�MJ(P A�P@� %�tV��2D�#b�y�%1i#M�7A�7��Y���'·�LK�ۻ�l�yv|�ｇ_L8>>f�&�ˬ��o����3H���_]+B݊�����v��y����cm�y��Mz�қ����u'�X,�N�|��G='�I���|���8??�֭[ܹs'��f�yNUU$��O?��Ç��_[{{��$��f�D�_���+S�����R�"���1�3KV&TJ�'���k�:�^ ��h����q��LK5�`MO�){CWꦧv%����H�(�b��&J�$[CT�����_����{�:��=�a��(4�жd:[ར��P�qDWUH�v�4`� a�� �@�0;=a����	]���!Ӄ�Tu�$/PJa���!d%�}�!PF#I����)q$q]K�S.m��#�N��ܽ�w~��g�[_G���-�$e^b�#d6F��� �=_��o1ڸ���U��(�1٫o�|{�v���_�'�&^q2.�����b5B���?��z	����.�^Y��/��O�<l-8��m��V
�u���T5y���wx�d�G)REk�t�5Q�eKS�(F�(�<��<\�>�����й{kם�Jκz[k�
�	!�J���EJ�'�X� �'Q����9:
ܪ�HB��_�3��i�!�@�݉���ǯ֚$������3\�}���Y�Fk�f���]f�s>��}���խ/A�s��~��OPڳ��t]�p0�H�,�@'1��خC-_�^��%�"�#Z�SwmH��Ӣ�"J3�Ԉʺ��=g���gT���k�JyRO�R���!�g{P�k�\���e����u�a:�����X�o%��d�JN�Y/��闻��'^�=��BI�� ��GxG3!8ím��gS�@�G��/Qv-eS�%�XÄ1��hb�ED��`N��@����U�L>��&(B_R���%q�A8�f���8M��dL-$.���ӳ)���g,f5��)��Rv.mr���<����h�=ۛW��g��k�뢘ڍ��m��6�A�n6`q�c>��"����W~��='
g��y =�	����ˊ[��k�D��J��*�Z��ٌ���\�as{����'HT�b�t�F�w2gZ='�rIV�g���ܸɍk������@�t�|Q�N�zK�Y�ڬ�2V�b�u|�W�]�QU��(������sNOO�y�&��۷�u�7n� $[[[�u��L�%�m����QJ����`0����<~�!o��6�����u]���ŧ�~���_��9;;����8N_������:�1	:�����_�W���?q)S�mO��ˆ�8�M9)��kZ�8Afe��qu{�,����w=�I�Lq(��g2��#f��aMPY��B���kQF�:�3	B�����>��ݿ���}���y���/�9��c�y#OE�Ej|Gm��a�<���]��Z��Qu5������D�a�Z6�`#����nLQ�2���&]C�5�����=��(�>���C�}vH'2�ؓ8O�c�k�t��M�FC6ӌ&$��
�0�r��IC$3揎��/�#��-�d��]���1�t���kT����5��!���e�~UH^6sy�KR����Uz�[bE([*�.����D "!>�g�$J�:ޕ,4�2����ײ�<���a�g�Sխ�E�HI��(Q�ܶ�löwí�F'@>���� p���	�;��r���IY�"YE�����L��i���=U�$;��B��{��}�Z�����lӴH2U��h�΄ �X��a����:3)!���L����!Qk��{Oc���)�4���M���e/�"l���=�`����e<.�Ic�c^,x��_ H/:��GX֗�ۊ��hW��02�[=�A?c���:�bY1�cʡÍ<n�K2ܦx������b�i+�U����d�"��&=��$!��T�"�@Ɉ^2"�N�C��T�"��H/�D�zZ���n�iCP�����~�ǌ�mN�#����b��ސ�(��Ǌ�+�EA"bF�	M&R<
���-RH[	H%�HJ���,!oXCٴT�4� c=�Y�����;�-!@�*#HU��mc��貦&�N#d�1�4*M1�s��g<<<�~�7qq̰��m�^k��=&�	˦aq*�Js�bʝ�(��f^������|�m%�R��2�+��9+k��7�1/�3]-y��O`^3��Ͽ�"y�tV�\���"d��-���mvtN�&�l�87�5Kz^����{z�&������ĭJF[��w�|;Gf#���>�B ��ۮ��Rb:�+�q,i�2�p�܈�Za���i[�sH%ɢ��ȓ�&.=ES�
As���9�~�5�f��p��R���C�s��G��GQ�5����T�E�8�ʕ��c�ɐ���zs�N�x������cΝ;�V��1/�c��ժ�ʕ�NOx��!'�GL�S�������dcģG�x�7xᅫܿ���7o��hC���Z��_�~�q�v�Q�RuBh�B�;�My�k�}b�pN��=Oyr����s��2�݌s[7h����aD�8e5;�b��>���.<U��Ti���=�p[��GD%6�0hh�lp�!P�s.���}d�7������}�ִ�������e�i[\k���rxx�1បMA�"2)9���'waUcIF#�o���ֆ<IY���*��ZL�8^���o�;��>���ʒ��n}�9q�<�Ӷ�~w�˩�_]�E�*�و֔�|�!���qN�@-Y�YE�O(W5y>DM&�._�|����	�/��ŕǷ����l|�1ʠl�5��ZH�� ����5�}-3��Ya�n�EH<+
"#(�
G�:!�
[�o�N�]��
�'#&����hi,m$�מ(��DE_[�˂Ţ��#�8�)IMKѴT�E�%�ڶd2e��H-q�ߒ��`���@CHS��0w�[�4f�\�d���H��ŶUHb�����4�\ʲ�VCk�gU��*ƹn<ꂒk82�G�>a%k�b��H��Q���e&tW���'�a����Eh<5+A���Cϳ�u�4�w,C)�u4��"�1���Lz�v69��1��l��	E��8G�8hGۖ�x��h@��,��� ۚ�y�Pw��c̺�:�܂m� ��H麹��<��Ͳ֒�������~��d2 �Q .J��R�c<��JM�B�`qĽ$�(J1��C�Q��"@u����Z8��:X���L�hmS���b�i&�;���8)C1�;d@�.�����UI��zy�;�Y�5��|������]��Q�$��k�F+I����c拂�|�0O���]�߽�4����۠��$u�h�
�^X|[3hI����8x�ʋ�����K������8f����*/+V��ܚ�c:��Rۍ.���QN%�,�K�|z̤ק)n�_>�D}��T%}���"�=�,�ـ�J.Rx��&�s���-!����ZK�B8�z�/)jK��DB�ZK�c�o?��bI�fx�X���$I(��sX�X���UQ�X,������yvwwё����uܹs��l�����^{�5<�GQ�����c��V+vwwIӔ_|���!/��駟2�L���`�s�=�1�{�)E�@J�+���`0�Ν;�L�iJ>3Ce=��w$�~�w~���^f5_�)k� h�~�����ξ�{"%���ST�����wBc˦de-a&�� �.�����Z#TL*S�R���US#����l�>����N�����:͙��t��j2��z�e^՚�tʽ����6�x��U���<���9�{�8�X-Y�4z����ܘ���ӌ�,�W��[ˍ�Oxn0 �c�4Cnl���i:�k�A	��/��y�0��b>;&�;`�d�)s��u5�|J~�<NKʲ!��ap�ɠ���7y��ߢ��l�(Mp}��	��⩌�Y���.��L/���,OI)����;�sxgqH�:Kme��%���,z�+ޕBz���Dz�N0R����7d9�:�غ��E4�
L0�Qu���yz#��QU+�HS�V�mM�d�2dD(RM�D�eEY�H)��$��ۆ,	�W��i��6%քF�i��ӏ�L&c��<Ii�E@��G�;w�ꊕ�t Ƌ������7��7���2x�O�A��Ҝ��>������a��ģ]�E��WX�E�A�dI�,�$Rk�y�!mZK��:���N�p�!��!��Ux�*�Y)u���VV˂�Ɉͭ	! Ó�}z�q��II%h��(@�y��5y?�gJ2O�n�t["p�:%�b���FD1�ɘb�R͏H�����A*b͒<Kj��1%%�٠-��L����8<�$�LN��
g,���~|�������MF�1��,���p||�1��X���1M��l�aY�E���K�e9������e�
4Dk)σ�9'��ĉ c���`>�����)���TOu�HO���:�^��H����C�+�l�1�#�g�ZK?�Qm��#��Ru�����A�G
�R��.�TE�ư,g,���T���!��Q-o�H#�/��&�4H��G=��|]��Ж���]R]�6aD�(��
�*t�.]�����{�����o�,\�~=�9>|����C>|��0�9>>�W�^E� �;::"MSv��f�;8�����`��~�����I�,�K>��3NOO���bkk��������s��}z���m�g6��9���#��߽��tΥф���osq�"'�s�vm%���RH���$��i�A�`�RT+uC�Ċ`~/�rw"�%ZJ,�ILݶ�MH��c���Y,��Ï��\�p�X�P(5�{l]������=����t�M���SKY�I�r����2�Ͱ����$��z%Qa�Q�h-9jVԍ�ɝ|x�g0��7����&�>�\�g<�������laM�����3����,R�p�)I���$b�I�I����Ɨ�r�Wj<${a������4O
���*�,#Cߦ$Z�`��FaI!�ru���-���?��}
��0�gk�~��i-C�CX�ݿ�.�5��� �%��z"S��h�%�#ʢ�*��4�\H���p0fZ5���z��v�=����F[�HGC��P��U�E����8$N:CkjBք��cj��DQD�k�
��&��f ��&Ob�4�&��$�'�Qۢ��M,QU�9��1�3��'���	��\c�#�:�Y��ERx�-����W��=��[�&���w(668],1.���q��؈MS�jV��K�W%ug����X	�i�%Z�X�q�D�;�y�Zi�Ԡ5u]�*�MI]E�\��5�,"�2�1E�j��Z���=�<�z��-��!�ш��1�b�E����^9Ϫ��������C/��iB���F E����^�!�^]�O�%�BRUa�@k�28V�~EAmy���0��N�|�;������������q��M��(W+f���)e�eyG�mKdI�9�k=mՒ&	
�I���q��#n���b�$�6�&lll����IW��`$$��K;#Qё--�h�R�lD��xGٴ�X!�����ɈӢ����P��mT��y�s��d��.Vθ��(�QB��ka@��
/d�0����<�x�JR��8Oy�����Ƀ��=~���,�Q�%eٹ�����:¹Ё���}��G��gv�Ʉ�,�����u�V06r�H�y�&J������F,>��#��7�N�쳱����c��>RJ<x@]����럲���s���։_���_�Ī�Z>��K��� t�0��ؾ���x��-Y�O����V�4�8K�"�T��T�A*M6�3�����>��%m�(J0N�c��>tC�cr?��H�w�=�9J[A_��S�� BE� uL�+N����~����o��H�0IG�^h����t���X�YLg�'%��$D��dQ�ko\���+�OBp��m��,Ky��1m�ppz���6
Iq�`+�`+�;�	[�[\���.����8=>d9/8],9�?�xz���-�l RR�*�1!�\�<�����V��A	M�u����4}�������3�[^���!;����߃Yt��g$d�)y�{���f`���Iޙ|�,p��B	�Y��#���pጲ#!��Z��ha������k�3-���������(�<�Q,K�G���m0)Z��ٌ���{�u���o���n3�CB�b4$����Z�BQ�!9��2����{�z���y�ˠ�HX�$�� P�c��`5]�%�c��<O0������L�p��z�^��i�vv}%�N	Ak-:(-�������S�S�ɂ���3���+n�x4�Nb&�J"�����okQk��a��U�~�8�R~����� ���'y�[�`ƭ��9�9�&c�+&����bE�4��a4`�`9[�#��60�>˓z��#��!�/^$�Y������iy\��,HJ�D��hK�ޓjM���f�>'��oVz�V �?�RBvz�4�F⼣?Pac�����ѣL��	��.2��\��ʡ�*kH���l�1-u�P%�V�͂T����j5�C�qUI��a���*T�
՜���ϱ�:�Hǘ�YKs�Q�RJ��9�Q��oQQF�9Q��h��N`��2�"�J
�������w~�����7��*�X�O��34��y�[���T���힋s�@I��AS�٬x��{�7n��Cd�I��<��V&���m`���Qｧ�k��#�9hE���l��w�w�z�*��c~��q�����P�9KQ,Bbc������%���jɃ+�*����<�֭[�9�)�HӜժ�ƍ�9�e]���/��֭[�n�m[��x�pzVk�����k����f�x��̖<޻�d��n���bDc�8T��̪����\�x#��F)����Q�����;wʯ(b�&T�2�8Ꚏ��j�dI:ء?q�����>����a3.^���4m�5%��ٖ��}�����f��kX	�I���kW����mZېnL��������ҕ�NO������C�ſ�C�<xğ�?����x4`����	H��Xq��Ü�t���'�S��t��h=Ҭˊb��k�1-��%M�ơ3����>i�3G۴��l�#�/�Ls���_�gV�?��aǆ���N��Z������Fl���j�m�u���t~,B���<[����-=y]���ޘ�Zp��b�ֹ�]����bM8�55�ф��	�q�qLY�=!������������?���q�c�m���c�:E�	ԍŶ�҈8�%��&y�sx�O]��ߪ
t�fض�b�C���)�Q�s��lN6H���p�k��ʥ��TIY-��A4��Xk��t��O|������\>2�0����VHW�˚'����y��e2�d���X���mN{[�uI����1X�q�ଡ�Z\�>�YD'��6茭3Xg�5A� kI�'���5��}���Y��4��b<����(��ff���`��2��{A?�^G9Y�R��o/#�)*�)��]������qRSC9/Q�)/���'���5e�]�G��,a��x��=K���C���0n5Q#�"Nc�eY�0�uG���m�i��{���w�����is6�[H)y��1�X0)&����"ȰNN�����!<ԗ5I�YV�4V��(뒺���mQB�9yϘf-?�Z�zdL.�
W8�MK;������|�H��f�,O�`��p���!��/��M2Ss��X���u�����g��g�JF��l��B�"��� �3�!$!֦F��aQ�ˇDQ��4�E�%E��JS6�,«�!8�PTU���>�CK�<e<�)�n���    IDATݢ55[[[���f�w� 	Z:�(��}l[��O���N4Q�%EQ2h�p�:W���3��?I����n��3M����
g`]4��$�����ѿ�g��$�'�[���[��P����]5XcH����������9ݧ���F����p��5R��A�u�i>�vΣ�
��>�7k�(A���� MJi��&�u�����8�/�3Ff��j���9�{§�~��/oaL�bU�(WHeS�Z��bVM͟��rtt�����(���f���'���7H�W߾Ƶ��Ai[�0%�"	ӓ=���a�Z�%\}�2Rx�'�G$Q��P��Z1����J�YN�(�#7-���oȏ�H�J�9��Е���K�|J��� @����G��%�{?��?A�C,�{�a!��g�O;��t�?z�����H��Q�8K��]1�Tձ�]>��#�>̺���ޑEnMU0����&��!<j0��=���ONH���V,N�FCP���}.x���KW�������������7��"�-��$IB�F,�C�g��j*L�t�G���u��L��9΅�&�b�6'��gkc����)�|�)Nkvϝ'.O8�O���H��H�����1�_�o�����=
� �����xo���K�	q1z����U���_���������	�ɐ��VM��	j�072HӔ�l��t���m[2�O)�%�����k\� E��.��L#�E	����VJ�	�Ci#�/�e9�	�8&RQ��V5mݰꒊ�ց@�Jj�i��;�� ���Kb���-RE�ۜkHz�Η�"���`����K�C���I�����1-���zc��8T��&�s�1�8�;,��h�h�&t�³���1��tJ���5͞�������kWy�ګ8�8<<��͛�~��κVppp�'��`4S?�G(\�tD�F�!JȮ �PB�%�A�|��&���ހ�P��KlkH�D�S-�l?w�w��=����'��R�6�~�|�"W�K�R*�|ِz�n�](��cE�ȿ*���`|��H�����z�:t�Jw邖X��xD�}�W_}7� ���Z�Ҙ�}�m>���|���|q���	uc�m0eI"��d�m�Ui�k����_���mNN���H���[o���o����<ǜ�Z���$��PI�d-�)���i:��(dY����"�y�w�D8 �<�m[�~j��6��f�u��ٿ��y*��!��7��'�L�\FKM�k,�s�T���(h��	��@c-Nz4a�����Y���c��b�ν.��|�0�EQ�"��do���mSq��(%x����6eU���#?~L]�`qt�n[�a�)�-�L���'S��$h6�}�O�Svww)�{��I��{���!�à��)N
�����:>LY�#�6��CڦĴ5�4��&4�P����Y�3���{�'���_a�fQ,�sMJ���T3z�6_�o3�?bh+v����\��������z��]����Y����(Uw���S�$�t�;���w"x�t�<�ΓMf��]�z):��������eK��)�X��B�Z�޾���e���;�޿����[��o�+�nA�,XU��Ucp^Q���љ[�i���H�|h��84\��.p��E6���L�S����F�)��/0����uĽ�z�t�4�ݳ�{��G��S�^�@K��Ax�V �G�l�1������$��w�6ΑE9��Gϧ$IĪ�x�4
���/�D<ass���'Oq��F�1��;�N�|�����p� ��i��DJ�f�aS
a���#]��+)���F2�L�{q�ţH�gB�gyp���jCGT��IM2�1�t�$IX=�G%�Ha���3���p��4b����'1ҁ�k��sf��U��px)0�b��u��hD���Ѣ$az<#�^��®PŒ�j H�x�y�Z�7�3#S7�A���(�5��T��|������/��ZK'�,�'H/Ϲz�*�^��W����!G�,�K���jU�>���}j
#���i"�aJ#/:���-=��U�@(���s��}^��2I�/�Ll���)�	�T�Sܨ�T1Ac��&$eYyv�B��Aj���lHrG�3�$J�ذ�t0p�[��eBop��J1�MqB�\�ʋWi�`4�)�q��iI��Hil[�d8��D�]0��{&�	/�pu=뭷�{)J).]��l6�'?��z���/�ꫡ({��>��k.^��ʕ+x/�}�6GGGDQļ˼�������{O��cww��h���^�.�loo�����8�B���e`���Z�u��9�����7_�7]�Z��g�+Z��R��zD���V��&���u�eEU�鱀	�U�{;_
)�z��i����ۅ�8s�s4�~�pT��O��MB]W�4��-ٿ������QT��S�L��~�t0`���"T֣2��7���o�Xl��p����h��_�����i889�?����V�9�������,�S�X �f��f�,��4���1��Iv&�8o�ɒ4�u�"��bE�ִ��El#��1ތP���aж�C��y�P��x�xf�%:�˳����ڟ]_����U���*��~M��;C�TǾ�;�X����Qk,�e=Ԏv�$��$S���K������7���m��p@?K�����s��y���ӟ��o�������׿ɕ�_��O>�����/n�fUդi����"Nr���xՍUگ�`�qD��g0̘�Ɯ?w��`�1�����C�'ǜ�ݤ�si���=�|t��U����/�إ#���"���ր�h�4I�yMS�]�b0�D��4UA�D�~��7H�\3?�K��E���UK.���x�
�=�b�"���d�ŗ�;���8w��'�i���y�bUc��H8|d>���X�A� hp�lL��w��xs�������%$i��=���x'-�~S��i�Uͩ)��t�G#[r$M�g62�{\�5n�1s�k�Z�i�dЧ�����Y��
ǩ2Tq�o�'sJ9%�,�H0.8z!5Ά�6�JZD�Yo�AG��.DD��![�}C��4F������.q�ʥK$Y��{�i�AD
�Y��j���w?���c�Tq����p��s���6��p���X	�����@��`��ޠ��"�ؖ�*zy��h��KxpD.43q����s�������q�[����?����J�d��p���U^��ߧH,�pA�5�����u�Сx�0gH�;K���Kuc� -z���p�u�:�4ZR5K�"�̠2GQ̹y�s��%e��Ĵ�~z�3�n�E��8 Q�(˂�>�)�N:c� ��x�">�a�D@0y�W�Z�����}�5��9�4����e�X��o��{��t:%���ı�x�s{ss��տ�G}ă�Ȳ�7�x���-��b<r��-QQ�q-�Z�
�vSJn�2���<:e0�����]��!BK����^ �YO�i��x�(��0��8o�Xİ������h���	��YU����c*�vI�)�Gl�����_���\�%���A��I�mjlQ��hH�899A+A�T��8R��>�|й.�l�����?�{ϻﾋiK��~�~?�O������V�u��A� �d������a��ł�bF�n�����틤*	Y�CZ�H��?<dUW�Ȣ���(�T%���HKo���i�A� �xn�<�Y�z��RƯ�
[������ub�����mAk��φ���`_#;&�0�2���=�%YY��3D�b��9
',�������
�$�R�s�����h0h�ZO�kT�����u&�o�}�*Kq�a^#�g�۠��Ű����*����e�x�d���}.��pxP����5o����:�Kݴ$��W��u���nݼ�g��Gwo1;=bY.)}E���QFaBc�ǶQ1���svv��<��,*��Sݿ�3-[[cr}��M�������'잿��t�<�8�`Ψ�B��6�^����""�!<6�rnS�!��I�S��C�x���#�Sc��I��K� &�&�d�ڛ_g�KDYΪu�H����Σ����sxx�������0ZΠ���Q�`F9�L����BG�$�G)��x��p�b��s
g��(I�BZ��(�
�$xf�E�7-2�G�$;����o~�C�r9��>J4ȶ���������%�4�h�Γ����i}Ki�x�! -d�>���"���x��F@mY�!�9�g�I��(J����F�-Jb�����	/^B��Gǡ�Lb櫂Y�"�S��ηy��KE�ݻw���g�e�iEX��8ʲ"MS�7���ZY*i0q�J߄Y��Ғ�1��&ۆ�!ᡗ��Ä�K�G�w��?�_9�CړS�?|�Z�99=B�.I�7��,y���=�2T�g3óMI�O�w??��E	]���g_sNf�mŕK}��>����YLKz�^x����_�%<@J�+��z����tg�a�t����/�ļ8��v��ڎ����.YQ�w����/�$I"vww���`�
��~�3�1�ʻﰽ�����[��g��hĵk����Y�}��ty�s��V�׮]c2	9�B��!���'ؚ��3������&��K���� �J o��E$:���(��T{	�$z>��5�p(����(T�%�e�bX���/�,e��`��h}�P �Ƕ5����E�1M��t�Ҷm@�@�y�B�R=�%[�ʆ�l�䓏���px�K�/0���ύ��E��d�m/:d�������^��uX�g��Q?���'�b��D��m�����c6����3VZ3�kN�!i<a�RJ5F��Gf������T�Nr^z�U�_{��O?������Y�h��:��v��K����9U>d�x�B��r@�6a:��U�ܜ�>�P�3�{x*-;�p����_�,��� |�4�\Ŕ�9�K���7��+�u����=���ͭ�?�����l������8:<�׾��\y��.g%�J�K_{��^{�f9eo�	����GOOY��óu�,���0�������ĉ�1��{�<�s���#"!������K�qz��'���4��w�r����������h6|8��
���)��It/'��ՠ�Kb욍�����`;I�I��x̋W^���W �4�^R��4�H�۴ԫ����'����=�?�!��)YSд+h�.A)�5
�C��:[kt�#���ŏ����"vFی��I�g��Y�qR���Y̧�M�����1}/X,K拂����*q�y�1�"�L�J2]-q�b'�T~��Fi|�R�JVeMދi�f6��;������]��ntg�`/�k�^"��6��$��/I����E���Ƅ���m�2�5u��>��s�y�w�4M��Ѵ5����f�eY0��*���	pf����lBam�~
��� ]����Ja��4JqV�\�X��4�#J%'�f�[Lےf	��	����?�}\�I��y���}���IO�����{�<���K��_�Y�3��k��c���Ō��/�[;X`1� �9�P\_�����=�]�]��M�JIʲ��@��tDk���(
666x��w�L&|��'ܾ}�8�R�|�u�B�y������\.���y��!/���Up��tC��)˒,��㰪��}�6����b�6�9�����1�(���ϲ���_�F�� �;�8w�������c�K����>�/b��|4
���5	K9�F��$���Ղ�\�kG�Dy�_V8٠u��Sƛ[��e6?�µx2��
�!J���\pkt&�AX���iI��4ɂYS��R�e�`1��e�1Н��؆8�0qL�̷�Ϳ��z>[���S.]�lP;Wu������7R��8gܘ���h%0>D��y�k����[T,�%�y���ﲽ�2�|�%T~�i{Don�ӄ�����o�C��zQ :�;/%V�.�H���Yq����S��/~�3"��gy��L]*�DT �:'�*�^�2X,�����z��Ĳwz���f|�"��i�aV�X�������c�|�-^�,fS�vw�1��'pr�Ϡ?�-N����'\�w�������K�(
v��'\~e��^ycCfD;=�B��$a����Wq��gkދ�3q6���8兗.��ք�~��߻��,e�Z%q��W���\������P��ŀ��<�m�$ �Y���^K��$�R)���C%�MG/]z��<��˂^�'�4��xƵW�Kԗ���(9��KR�o�lE_�X�ǹ:���/�^#�F�'D���7�dg�"�Ҙ�2`,B�;c��S�OY,g���lGV5��);�F6�F��F�؂��xԶ,��9�X%�D��j��VJN���W8"D��:M�z�v�I���wn]��SBwDg��\,
��jQF˺`�Z���׿�2�_��d�N�����ɓ'ܻ}�4��{=z,a�a>���a�_�%����/?��ͬv(����4N�R�V4mI]-�B�&���)�U��[O;]Һ���Y �D2"��.PZ3MPu��Ƅ|8舆-V��4�TD|�;������L����=�]�2s�Hy��o����]<�+��]����[_0��?%�m.�Tn�s;����Yv�y(�&<'�2�4��7�0Ԅ��%�/?�T�T?�C����h���t΍Bj������t-eY"�d{{�o~��c�_��g�}�M����1��Or]���,wɽ�P � .�(J��m�ew��ݫ�=33�|�鉙qD�������l˲H����J,�^��]�2��D�1�(���y�y��>����N�C��\�z����%)�sf����M�]�������T@tFɯ(����ѣGE�,��ɄW_}��/.O�q8��s{������=��S�Z���N�< ��Y-��dq�A�����s��-6����1=�c6�$��Y3+,�La��#/*�+�}M7]ź�aY��'$�q�"MS�H/�ҘR���:�����6�MGO��b���)r2�����:O&غFᩫ������&��\@Jɝ;�B�Q����6�/�ȇ~��ppp�x4BIIEX���b��K�C��E���|:E8PRb8,�RH�*�5Q�غ�+ͅWnp���tё��P��ѐ4QĽ�� !;�C��s�,!DCr�K����������nQp�o1�v�Yÿ���b��D2�8�|���|S�7��V][r�������M��9�v�|Zpr����X��d�y���^���(�#^y�m�/�ȧ���'����⫛r��1[�/r��+����]�i�k��T�V�CUQEx�L������Ib�j���1�%��\��˗�)�>bv�}I��-Q�Pec��k���a�F��Ra9��}묣�̘%>RD&�M�.���b榢%,q"�,$��.\B )ʒV��D⫚n���r�S��QIJm���-�����Tu�}G8�zr[�:߈�NQ 0gX�[�|�.\�������"���u��J�"f�n�մb>9C,�{3.薚pFQׂ���"��Ŝ��ڔt}�����E�5VF ���6�z���d�����\.�_���zޟ��ߋ7��52�t�-�8bg��_���/���%J�(^�����F`�ct6^&��yN]�R�ISz���zm�|>H���ok�N5緷�qrv�� �oБ���'DiB�ա7�t��1�j/@y�EAUIV����B�M�J��b���I��˯�[�?"��@6�I&%nrL���Z�������jJ�f�w�~��lQ�6������ڌ_�16,O��M1p �I�&	���t�:�Mɪ�k�n����6�_x�?��?�>`6���Ӳ\���,ј���Z��3�]��[o��֚�>���?��(���z��	^�8M8���������Wo���	�v��|�;h��}�6��n�����
#��|�!�v:�.�����cn߾����~�~?��Ӵ(��b�s"-Rt�����������	���8�R�V�E�E�1�� x�?=��밹��6�    IDATF/!i��X�l�h<�w/p8������}�lĎ��V*�����M'ċ�Ӥy6I(�F'1�� �tK��ݭ.I����Ez�.Y�1��{����!�,c������G8k�$1��c�����q���,�(˒[7o�}���yI;|��_�ּt��|���++kıF���N�G���	d?Q�F�����Alh}��.g�����/|�[T�S?���_~�y<�*A�oQ������ti���)���ry/�C����g#_����Ιl���Ͳ w�z�����mF�W����0�ɜ%E��`�)�צ�m�֚���#f��w�{���ֿO�� �S�[W7�������3�ߧ��9==�l�t���[��ӄV�Og�O��&V��fU \���>urDUUlllp��"I8z����>�A����}��+��}��.zxF7����G�^�i@Շt̠�|vU�]����}h�J�D(�8ąC֒��_���c֯��::F�1��Q��#V���E�덠�4�P�v��1:G��tYU{;��TEN]D�Zi��AtЀ���/��xO�,u�l^���)���^[d�4��*�$�-���|6��,C:C5�¼ħ^J�N�Y��k����
Ó;���q�$������o���Gԋ)g#��������}:��b���L���AΉ`)���|<P �8jkh��ٌ|t��k�����U
a@i0u��5�(�����Sf�)Q���0^X]]��UC��8:9�s�l�����u�g'CΝ��ښ'O�P�:i�3Z*�^�@�ߢ25.�T�X@�(�G(���ZA1��wx�xfy���#�����rV&\|�:��&S7E�v���w�wo�^x�K����\�DQgĭ�ސ{?~�G�JK)�sZ)$�d%��->��V���\d� r����.���m�.�X���|��ʀv��N�%/@��yN����1&jR�:(-������+��\�����m����,�BMk<x���1�{�\��R���C��͆�������z��g?`gg���a�X�(�~,�:��^��`Bo��θq��Ʉ�d�J�5���V �����.��ߤ67�F�~�t>G�t�r�TZ�f�Z�F@Ƿ��x||ʤ3hEt5$*A!���FR�u��V�Vf�eY`eC$kDJUU��x����!V$�6��c�UiXY�r��K�x�4n�Q�����իW����?��ʹ�-����#��t�x$�<'�����F	+���X�^���ʓ��R�Z-���7��Y Y�T�4j�(�JG���)�$h=�$"m'�Z��ǿ�?�nt��2>�O�����r9Z!�5��`l����/"C��6b:/�Vx����O����떟�9Q^�c�����8B�ָ��~3�4Im`k�W�W�h�7�s�4����������7��\&��R�錼4H���;�`k��~F�I����A{�׾�[\�u=dxvB�g�m1������p�N�bO�53/(Ua��\�ܹs�Zm���۷(f�I���ֱ��ʫ�/Ү����o8��3��P��q;���n,�a���K��)���~w���|h��E;_)4�X������}6�A��S�8A疸.&���2>;����֊���xvJ>��LE�IH;1Q+�����㓧�.G��	:��j�S�F�ݬ.�|1%�D�XPU9�d�|�016/1��/!j��Mw$[]��ed�c��QL�S��:�w���v������O^��{��/]������8�V)*TI���-�|8�2�w��vD,e�T�:Ո
�ٲ��(Tk��	JFA��=Z
����Ni�&\Z[o�2G�1J�N��,o��I�CyCڊ��'�QJ���$�qqL�D|y�.�����T�f:����Q���G���8;�Q���v�urS�p�����O6m+k��m��0�O&ت��.u;�(bD�K4���n��!q5e���Ӛ>%���x���_��9{?{����a���7+�.�/`by*����s�E���k!�M�K/��}�p0�H���~ ���.������=:�.�^/�[��CG�YteP������(��,6�8\�ũ�7��fee�W^y%�!�<|��=�ϟ�ܹs���+c888b8�R����I[A����+D�8.Z�.\�ʕ+lllP����"��]'Z��QBЉb�o���]ǘ�7��=�5<��OhiI�k�k��V*]�q&'MI+%�. �#�Z�C��0�{J�9+3"WK�$�#����챵1�֡�d<�~�s)q�B�{$*eug������_$J�l��&I"�Xb�EHI�j�Mg\��lop�����p�i"����_���㝥�b�iG�4�<��rVz}�����(;�t��.e��)JK��	D"h���AVfD1���:���>���ɐ�j]��.в��d�*���ß���&��]zZa�u�-��5�/�v�#�[�v�<�w�ܜ
W8�I^"�G�����C��J�\�(�n��`P��I��NQ!?��ZA�\��\���spp����%~�Ο���]���o��.��
�� A�׸p}�g��c�_���wɲ��,�*���0��"bI�������jwy��1}�	���\��0�k6ϯ�����
���_��ݿ�5�It���D� �5���2� ��8���|uo���
�%t� '| "96XA�)e9�[�N�(��ziHkC��>���[��ھL�t�e�k�O��v^��DQ|�z^����ㇴkCG̽#�Ԙ�B�
g"��i7�?)QJ����ݿ�Õ6���6�ZF�G�+�z�<u���Z�ݔ��D���8�PM��l��f���HDGSaӍ��%B��s�m^�7��ڕ̾����Ԁ��ר67���7��{����È����w�@ٴ-��LJ�s��o$2,҃NR�҈J��"�c�ZR!��p�O�Q�s_`8�3�8��c>:%�F�V��ʀ�~���\�|�V�"�cV���}:�M踠Vq� �E��!T�|7N0��n���ft�.� ��G"�9<<${�ǩ1ȭ9���i55W/_acVr�������d��.u��QYA�GDV`2�f����"��1i\P���d�{m���_�#��Gl���gAh�P5��!�{�W$�=^����/��l2��}�U�"��.3�v�?�����98<���n�Ե
��\
0Ue�ȣ��`m͝�����`X�K��bc��D@���?�ɓ'�9::Z���ݻ�d2Z*����=Opm28�<�C�p#��N����)�|�	���!��>Y������O/��xvm����?}�/����G���������F1�٘��kyO���F=�tM�Ą$B�[���R0�ft��*�О���I��`�DkI� ���C�-��g,V8�|��k�Q¹sy㻿�΋�1����Q��Ca����f���\�>����������hXy ��u�QE�s��#U���I��BxAmJ�<��Jɲ`�L���`@�nQ��F8Q5��`e�)F8|�B��X�NU@��3s5炈���[ﲙ���Cq�.z���`�![/�C]=G�f���,߸����������m�k��}b�\3W�E@��.PDU��C��y���oZ��>�>�J
YPVSV���1�Ͽ���A��`��F7�ŃG)�	�o}����y�������-u���4i�Fv�VƔYI>ͩ��퐊%t,n�/Q~�ã>��6Ov���3���)��x��W_筷�`��9~�>��,c�#�P�+�ܐ&�,R�&�N.�/_-~�D���iSI��!�7�	mn%��eR�X��A*��E!�"��g�5� vw9�.�}8�1�`��CYS���^%`+�O&G*4$r! r,�:��%�bL��$dy��p�����@h��t��0�B�#�
�%���oI����y�p9�ռ����SqVK6�>y2�x�eV��H6q�o�����T	ꥷx���|�m��� �����#�eN-"�5JX�@�7��^����o�-��"�Q؂4��V3���t�k-��]�û7��j��铯Ȋ)E5�#@Ǵ��_����}^��2UQbˊk���%�̫��x�fܡ��R��#���t(���L:}��YM��T�2ܽC5�qy�}z�;:bVV�n��V���w�w�vS��\ȧ��s��L/N)m�j4B�eȍ���^x�J��l>a��"��z�/�*�����c��>��$�Z@�P�LAKkj���=���m� �fY�����gI玳�Y]]gG{5�s��b�ּp�����_RW*ҍ�F��ڄv�1U��P5�JG�R�� eY� �&���8��`y�O����ï��~�芪i�*���K�\�,2 Z�'''|*lJu��u�撠罥,���l�pL-�6˲d��ÿ����+9��N��I��;L~/��.Z�A��I��%4Rh��0��D:\lY�c�*cs�Ɍ���}E�E�,������^�d-Q'
Ib+�y���4���Uνx��Ή�B�t$d��2fv6���c�����^#�������C~�����*�
�r���l]1�GTU�4_X��JqF��6R�β��2�:�pUQ�DDxRDK�W���NW�J#l��1��l�)+�q���_�;������I�q��������Or��C^z�{+]�o}�R��J0P/��" Լ���l��I�|�X�����{�Q�[Ե0��
�S��b�a R�:���&��zK-!�����J
4o>�DF�����HA5�~�.[{����Ѝ�>�� ���.�{�L�>��1�?���W^���7��؂HC�ѢZ�rA����(��V�E;iR��L�9�}���._�?a4���Z'e4��Em�z�U���������w~����n��Z���O-�l�atx<ZI�gJEH��$1�����zQ5��L��<W��Fh��$vN=>AۂY1'k'���ߢ��p�v6D
I"BEl�[W$�c��2��5�_�ehwyI^[�*�D�I"b[���T�A���9�l��zCe@[0��BE8���
�=ڋB��)FD8g�J��]�кa�W1y��R}����tDLy6��sV7�`
�)YG�GUԔE���.�o���o�6;�����^�"�m ����T�J,����	��F��V2��q��4uT�1:q�6χ�
�W9��>
W�*Pi�JUT�a�
Y�̊������v��7��������!�x�Q�1��9h�+I��(�"8�󌕕D�����2/p���`�YD^��
�4M)Ƨ�\h��� =J���
qg�{]�"�Ԕ��m�(�E	ǶF�6����q�7�5U^a;)�|�Њ�����\!��1��������#��xe�-?��IIU�υA��.d( �8
\g��#$^:�>���>�CZE��`S��$��߼�8���[d��P�h����� f-�_��\6�/	�a�"�QJI�g�}+d7�*0��B;�H��yh-��z�`�ѡ#��[ڸ��~���K��9�z�4^�[�Y� C,���pH����쀸��I����W��޺ER�`J����7"�pZt��^d�8防r�EM��gh��v��|<�ٚn��R1���GST�4�ט�f��Ǖ5�Z]�T)�.^�_â���{A���.��O��'�p||�J5��
��g���a2AՆ��;Y�P{Ls�A#���A&�.���FM״?X�;M��H���n����:i#�Y�H-�Nk���jK�=�5hk�8�D��fT�\��|���(<`��Y��^�q��^����s2!N���2�S�ʠ� FAGa��)t�>Ѹ�\325� / �Y�b�=�E��� s/���L��8xu�	�q7��2U8�+�h���K@��:�,���Ŷ��������/�����Xc��A���p��h��������p�/_}���sHS{K'M����<GzOn
���~:��}��S�s����$�8��Dq~p��s\�q�����or���b��mV�hyo�X�D�7y>�p�l:`�Y�DJ�TϮկ{h�,B��k�˓Sxfi�A9���@�1饫��?]"Mc*]����k��6(<S3�.+�"���`��,�[u]#+KQd8U#&��?��٣���b:y�1��(��/�nn "��L�?�#z�:�>���-�6B�3��(���Gk͠nQ�6��!:k�Ce%����(�)��^�������+��~��>~5��\z���-2��g^�O�ᔢ}kӜ$��zRV��I;��Ւ��k�}�ll��4�
+j|�q|i�t̅g^���1.��󊲘q6qZ���㏨����qe��SVP���&����t��JǼ-i]�d^��f��� +��,�H�iQ�������t��!C��!tD9������N�,2ј~�du.�c��������G��o���w�v�!�@:��Y�s#bUQG�Wt������A���c�H������p�CVx��<�5�H��a�g�H77�{딓��d��qL%-�����
S�h%��O�!d�s�rc��/���Ο?�]YP�(�(
�,k6�`WI[A���Y�>dY(ƪ�
�p6�N�CY���EX�r߯���o#B<���Dc��Cq�����������V,�;�vUr�ע��G��6��baF�H'UP TDQfL�a0�`�b��Q�t�&JS��1�|Q��)��P:!U)Z��^K��%3����|F;�AFH�(ꊙ�X��`Vdqt���![J��v����l�l��G��8D�:��̐q�5[״dh�[!�J�k�A�������6/^�N��ӣ!O�w)�"t=�6��k���M��sw��l�ۭt����i�F8G�_e����u�����y�_�+��O�ՖK��}���}��9�x��s�?b���Z-����%D��F>�QW����<W��w7�ş�րC(���L������R�w1B�����MU��o0�!����HD���(LA9;c5��[-��V�물��h>���Gd�G��2���S����iwt�=�&+0y	�१rɫ�"Q1v:#^��"�l�Ղ��&��Z��;/s�K�������ݟ�qp��;b!)l�� �Dx����-�k*=�&��/Fi���F/Ă���B���#H����bQ�O"cDY���$i�j%T��B;��r%5
��M(&��x� �0�&�n!��*��C"To����Ls��!�Y���I�`�+?��l��7�6�����/x��;/^&w5Mc<�:=�����G�&�Q4�+B
'pVQ%�K��e�I��`���6��ul�6��e�~�0��9��3�����o�������{�^�����ҳB��-�Dj*f�q��V)�o����5A3	�T�@mI�F�KX|M^�f��3��9:9��V�Q�k��
��e�������ұ	����6�ֿ��$��<�I�(���I����
�Ut��&4fck�V�EYې���M�H��V�v�K�,�	;L���?� ���5Z�Z���U|�Ú�֤�:>�0��ɌhU7��!nїi6��9ВkԼ�l>
��2��`a�>��s�n|��W�cV֙�*���pt}:q����v�R���x�)�����MY��b-�>��]�v����0ư���͛7��/�tUUp�����dgg�Mloo�������0�����K���fs6loo����R���� �t�q��2�{���.+++���/�[Y��A %�A�B��f�Z-�T���뼴s�2���?!�ߧ�O�kK�����,�~�`�-��2<�Ե`^X�.l�	��;�QJ�Ɉ��	REH<�)�����C*�X�E̫	�)��W̟�']['7��dL��E��?�g��$;=����������5j:!��x6��,U*�V����M�5i��H��}AA��$ed-����ǿ�i1E>y��<?�Z�    IDAT���Ǐ�L���a���`���ee}�����?|L~�.b:#��`3�����R�lm�����g�f 5��	�R���c�����UA]���5!3n��RJ#�Yf�{�LDLCF�����u.������E����&1��'��\c��_I�
-$Z�M~�a�B"�����!��d	=m9��}��#6^���6cѠ�7_{�Qg��Ov��1�v������R��%1g��V�8��!u�9��ϱ��
gk�$�V�o�s�E6��ď�p���'�;ڣ�I�I���e��y�>�ǑF����%��H���"�"���e��'�JM8OUL0�w��'�Z�@����D��(�@/Z�@r5�EK�wH4?H�(��ģk�1�|�cGg�U�Ob�Tho�i�D�I#q���ј��������ID$��)m�ùMG`ms�#T�J"tJ��Q�೚~+B` a@���3�ftv����cz�?�W���JG���/^�������R
ur���C�t��N���]�Q<W�.��3x�)�)�W����g��B�Y�b�@h٠���&��NB��S+���6:v��$ni�`Z�UNm-^x���HJr⽔(��}6�/��<�t4%5�8A	IU[���8�25���J�����>�~%XI�[�C˄����!7[V����0's����GFm<QK"��:�p�d$�Dג�@�#�'��e"��@o\��:�D�SQ�E#�i�]�| �GX�� �PB6�"�p
mzTU̓aάv$�U�V��gr�+L��Oǔ�R���)�>`+B�|v��y�Ç�M�\�r��t���)Y�q��y�^����	�n��^{�,+V�~�U?~�o�����l��F����K���ܿ�G����x�7�9����8gȲ���{._�L���޽{ ������쐦)O�����#�����@Ol�BGtW�y�M���D�3�����]v�cZI�Œ>(�D�!aA`��6�`7U*�K8��}�@Q�0�%�tFUT8ch�9y@��g�|N5�0���r�O@�he��=e���n�J����CQTV9�����rt�n P�A����(E-���jd-�|Q(ڭ��:\�b����luf����Ͼ���TG�R��
%b�(!?N�nm�:B�hR'�5�C�ʣځiR���e�v���tksa�i]1.N��%����O~��û ��Ԡ��Ϝ������&k�A#���������" ��"|������i�����Mؓ���(�ä�xg;�[vKY�����l4��K��2�NI������̰��Cg��)�N�����&cF����v�w��$'�+T��emѽ>�+:i���;�/����z��j+b|�#��>�wF:>a�ۥВYz�
!�D.�@Q��xg����/��y��֌�սpx,�.B?'�EK3@1�R������/|�����T�Z�¡��&�SiP[��qCB
m����QXW�O�X��ZC=����XY�1%���3������Aq|p¹�y�����[�(�v�(Ex���=e=gby����?� �S��XK�l���OI��R���{\�r��/"�e]A-(��1��<e�~����/h�3T��LN�ty=�1B�E�HW�b��G<��9��6���4�(�� e�6���$�I1U�ȳ���J-,EQP�%�"'�𘼤�Ͱ���K�0��q���;�2Ҵ�+�rij��B��gԽ.$1�f�e��@D1Q+E�z��o=^EH������,S�'����"���:�p�)f����*$��Eb+&՜
�0I1�AH��XᰮFzq0��3e*M��<�C�6��~�Bv�HT�p��HEh������I���3�ϱ6�c��)E�Ĳ=����un��޽{������ΣG��s� ��� |��g�u��˗����,��O������˗/��_P7^}�._l���3����s�?���,y�7����Ν;ܺu��l�7��M�qp�G��r��6~���W�\��ŋdY��و$������O����'���gl\��|�[l\��?@�WdH����٩D4Q�B�E
t+�5]�y���3>�b�C����k��iԬ7J��^;B`�Js���O���|�����%�jZ�6=�G�O�0�L����+���3N����э}jV�H�XM�.�iM�uUQE)
gpUA,=>�%u�ΐ�DxCV�TJ0�	*邮(&�P�E���F-*E;���A�o�-��XR����r��x������ē{��2�(�6��z�5��tHup�\p�i��8Y��.�]c�t��ryz_�������'e�G���d��&q�J��F����/��퐍���8A�ăgU�F���v<#btm�#���Ɔ�=N��A����W�{���UIn
�ќ��(�2�[�C	OL��mZ(�\����s���.ٽ����O�}���0������%����|��҃�L(����kE�!{⡽�H�N�p��.�C�?��e�LJl����fԜ:�o��-�d�z����p�)|�B�]h�.�������/�΅
�����k�R�Z"�N�P��a���):vHW�?���K_d��R��<�P8C�l�h.�P5���R��"J2MQN"�b^N�*V��b�{�������{ȁF9G:���<; >�������o1>=c>��j+	�����.I��4�uTyF�QB+�2�T�'��ƴ-j*�i(����F�Q�X#����U�lb �|e�pTe��+"�	�[�"���u�U��R�N���O:��dg	�e�{����;�8������� ��M���th�)"�qq@�
kpe��:ziB$�$��0�2:Q��RL�}Z+mF�1�f7�[���`���"l��X�� <$J"����{�y�s!	�{��qS蚠^��Mw2)��i��MHj�n���+F�5�7�u��c*��<�����0o:�A#���v����߸q�/�����}&�I�H4���x�$ͭ1�Y�X��ի�y�t:�n��p�{����)o��fj�L���I���C��1���8o8<���㇁���kh�)��n������e�+�^��d� ��'9=����Y8�.:��:/	���F�KX����N �;-TQڊ���u��H<e���*�L��,:�qᵷ�;b����s0��R*@,�9|>��|aCH�ɉ�l2���ۜk��[]|�pRQ���V��~��耞R���j�Y}훰�FQ�h���i�I���V�VB�N(�b6Ǩ�n7��ߴ͵�P�J�2�4�r�et��
�+�qBb�g������-ֿ�J\h
�9�(�!X{�m�/s�;�����?�*$�@x6��u�8aD`h,X+�a��7�}�����(/�������y����"r�峬��0d����e�(:�mB��xv���B8M�,�s8�Qi�h��kC_u)�g�|tL|�>��&��$/�t4S�[�j�,��Aw@�
x�C�Y$=]��UE�z�+�x�2�����;����m����A�QH��1���9J):�����o��i�;�q"�-
���y���8x�-�_���M�F����=�s����%콞-��;��
;�ts�F�@ 	RRbP�biF#�������p��/~��eW�l�eY5���#iH��Dj�x���O�q?���=@��b�}y�>������o@'c-U]�3j�-O�+����	@<�5F��J�◴&�n�ua&�TbMYWh���[j�H"�%R{t�P$�i��cmC�H�@����x��l�~���x�����²X,P2�1�as���f�P��"cFN�=���,~P 3˻wߤ���[o��]��?��h�0HzTT�,v�A]��4�,�T�A��K��?�F7/��M�����i%������5����`���,h\�m�"��j&���1eE�/(�����Z�3��]*m��C�[kz�:�ID��@:��
-��-�$��Q"���(+"�HX,f8fؐz	�A*���a���r:e�װqN3/���C�,a7�qA�`��\{�*O~����;<FR��`*FI���@Eqh��5�[����U��Ȑ t����e7K�9�Be,z���~M�ST��90�%���E�LR�i(G�Z����� y���8���&Ukx�Q�>��#����g�������c2�`�Y"����B ������^������oq��%�6wZZ_h�_�v��~��A5n��U��n�1���c�՟��:,��ri��	��y���;����/��y��������~�z|B_;�Ё����!�l�	-`K�'Ako�ʚHxJaLM1�B:L��»p������'lZ���ϿB�8fqx��W^DF1��d=�(�Ai���W�ݒܔ8%�Ƨ��W�y��`��lX`p�c�z̓]�՘�T"Fo^��7���W_c��؊X9��B*�������D-;I"-�"M�%Dm2��B�Ľcf�Sd���1��u1T��ɔ��.Y��."2!I�z5� "��P&fg�"�l����	��=ִR��V�T�|��ڇ�z8�[B��{��O�D��I���Z�[�~H�����O׶��?�O#<K#$u7�n}��X��*AyIe���I~J,cT�0k,�VӠ����>��	������=�o�D�?��ŋd�}�$e8ᅧ�
�k&���w���oQ]����t6g|�>��#�U� �Hk���D��׋��� �g�-�-���H�:pʣ�X��t�9]��L��`�Æ���.�%���8뉥Wcꠓ)�/J���G��{k@
d�p�)�n.y�B��k���oB��x�ZR��=H�TH�if3"!�mg &p`���������F)�'T��Z��]�����5!(�9���G�J���hOO+\��yI�k�ї#^�ʷy�_�	����#�ه���i�+" V��P�9+�1w���G�ǳ�/�
�ϧ�(C��?�6�K�Q��7�n��⌣*J�E�������تF���OiLE����sv��/(N��%ɵ�����KeL�%q�9$�H3�C{)N�Ak8ֽ�$IH��ʪB7	C�%��dsD,*���G<��;D~�����g���p�`���?�c.<w����ܽ�����!�8z���b�/�@_�B�bQ6OK~,�H�l�3�-߶�KCӷ9Qi9YT�6v�T��7�����Q���:�T}-����9�T���c�r^/�������2�ei/��?��>s�W_}��>���b�|>�Z�h4�(
�1�D�A�s7_�ҥK�D�ѣ��d�?�)�?�<W�^�'?�	�Ν���kL&v��Y0�i\`�Mo�'N�%��r��.�RN���������\�2~t��H��$Ⱥ��IR���6t�TΉ����ޑ��bt�P�s�/��UH-@I�lB�6H�β����'��WΠ���P��'{��{���-�҈�^�᭣�'����t�</�![�����~��c�	:��W��W�xR�Ò��dD�gv�j�>�KW��A+�U5�Lh�U�8�	G#k�������&���{��b9��I����q��U���vFZ&w����b���pz�'����;�׷��^v�,��)~1Gi�O���r'$~��H_�8O��D=�LZ��=ۖ������Ԕ*b�,R%B`�tH|�RaX,r��Z�n�9�ЧXQI,4ySSS���Xd$�>Ʃ�볱�!�Ţ �����D)h��2�Qk�������f[�OP�l��|L�{@��H)�i���y懛<Q����!�N��bM���C��K��cN��&�n�����	eQc]�$�
mԀ�����jKj�ѓ\&�DI��E�$�B�Z5������g���UK����2�C�?wgH�p�=M�X��Xi���%m��������zAK�o���r�� R ��(O��m�v��>o�L��+�:�B��Z�sr%�3Xk-��LH���P5Q)��	IoH�OP�-���F|n�+F�/s���M� ީ���*�,t챥'�g�H����ף,�A%�X@<_J�&q��EM�T!(T���|����;G]7%7o�5��,Ǹ�5�C�kj��܏�4Qɬ�TB�D"�g���p��mE8Oc;Nv\Քd Gkk$I����� �8�rA�)R-���H�)��5���W��/�ė��_1��A�0ϏI�u*s��/r��W����9e|����w���o�*�׶�<��>襎���'�R���#n>���k��Dq��,��W_G6����>�|�joI��UJTOg�{н�R���\�|��z�����y��W�t�u�\[kɲ�������������dY����rk�ϲ~)�t�������������+W�E���[&6կ���c0m��b�L���}�0�5i��{p@T�F�S�
GT9*�!�Ŋ}p��UMԪFJ)����R�pZa4��P:$5�#��� �	E^���L�~ȿ���[D/C���`^�Y��T�)B�s�ơ�
�a�3|�OgL�){�f$QJ�B��D?����ˀ1-�t1���w���o�#hG"F�h�g�D��ek���ـ8�A�s,N�A0O�c,	Q���i-����8ez�}�j<�b�!�%����T�£f���J2H��cQ�H�/�@G�$ђ���s�b��P������n�'�����G	�0!j����a��9JFK�� !z�*�^RIH�_W��#ED�em$�2�I��n:����,�V$��9�Q��EO����H��n���-��cd�z�in:�|r���=��e�iS4�ƒhM��l�h8�#�QL?JX�Pk`���!$��pf��×�u�sp��/)��!t��9�f�q5��eWr�5�Cm\DuZ��D��SZ�������	��k��	� !�KdG� ���n=x�G��nV.&?���*j���,_��/�*���u����=�l��_�L��G_�h+��9BXFCM�u��6%��$qB6Z��Fk��N�F��]�q�-H-i��
����zt�Fo�O�D�Ǽ���0{p��6H�R��[74Qн.�S�x�`���C� �d�/h��B��75nV�Ɉ��P����g?c��^A�PZ��2�F�(H�갱�!��5�����#��H��O��rU�}D�̦%��
Elnm�J��9�*�L(�s4�)�'����>N���뛛̏y����)���-�������Z�g��{N~j��w蟿���8�$��G?�qZF��b���k;��(�q�rS���rE>d>������w�}�o�������c�^����_���i�f�y��9w��eoo��`���}��1J)._���/�LY���c>|�R�,˘L&K��b�b���W^��ի��{��tID��������n>���飏��������9�W����A��cCt<*[���8��A*G�#Q��[���X�xKmkb�Ph��	f>G�Fz�V���5�z��Rn0l[�U]S��!%d�>&�Li��!�9�|LiJXkȧc�����ЅcV�ڡ�cS)|_3�Jz�B(8<>��"d������K/Ǣg�N�}����.WJB(�i�Y�Q9%�ˊ�t�}q�r�!,u�ceB�DA�s�Q�����R�i�x�&g�� ��G7��45��
U��H%�և�؂჈�Q��9�%�ʊ6�[6O����9�c2�
��
�u%V�7�ĜK�1��^4���u�M��:�	�����(#�i����V����Y�q�ʔA�I�g mӠ�g]+����qJ�֋)1� 
_-�a/�*(h��r>c|p�����G���ĮVǹ��I���샱�w"�o9C]U�uپ^!��;��.�u�z�J���X��qf#H
;E=�fƾ��u�d[�)aY�J�(N������y�_��Y�ᓔ�O�{ed�T�=��ʵ���wRh-u$���1<Lf|    IDAT�������hې�}���<��b+�V����JѵeM�̭	�B��'꾤%pNPUu ��k<��d����~��?$ٸt�<0�sD,��d<9!���l���H!�����◒��0xL�7]9��iuM/M�"M"<N&�c�<�$�0��/C��
�t��� �8i�܃�NR�,%�S�d"!���g��׷��������+��1��#�f��/?��׾���Oz�`��#���d���������n�^�j~Ł���O�m-��+x�O����z���L�j�ͧ4q�X�ܩ�Ǔ'x�ɢh�X�������jba���*>|�+MI���|�[o�պ�����szz�;������bY�w�n����;,?�ܸq!������������Cf��R'�L�������'�c�{�=��f�d�����Zé��w�}�����|�gx�/�ѽ��ctԃ%�3xtv���)-�b�Q|hg'4�X�]�t��TDQ��]��,��=�s���y4���/�?�Okk����TDJ�4Ͳ�px�4!��=!?9��J��qq�g-��ɔyY�x�n�:�T���On�=���[N
��ָ���]��
eUgq�ķ�>hj�	t��VqD��ڃ=xc�qL�@�A�8r�d)��������=vC�;��r�x=�aP�ufӂ���Z�
�����%d1�-j����TBR$��Ӕ�6T�����
���ؖq �
Oi-������[��l�%��D�f�!"c�x��SZ�0֍��k�,ySЏ%#��F�M;��cd��e�
fiM�� ��f-#E�qpW�TG�	F
�$.����'-z��B��X���Y;z�$�T�M�� V͛�Mr�>g�tD+^%����XF�v���H/ׯkײ1����H�Z�O�<]�_=�$���8����lA�QG���!�Dk�O��e�'-B�n�ס
�
��� ~�Z�w-��{�[A���7�b��=ӂ��
;t�?FYYj穑�:�Y�Y�q'����X��Ћ�x��K�� h�@U��֥�(�8��
"���zK"<���4j��n�����p�
��M��89=�9(kk��TU�l2a>�����k�D�p>�������)��ZlY��� g���Tx^i��G�qD�$	I�`	�|�$�RT� U�Jjx3�3s%�l�����;l<s���]�7�"�����]6|C�w�����W��ٯ�&GMAUhdܐ��������_YKq<f�4���%��1�ܲZ�gs�O;ى�����f��E<��42bQ,�\;Ǖk����r��HШDQZh�í c���.�]�;BG��_��< 
[��x:a��d�T�eB��f�UU1����^�x<孷~��[I���'c��>��?����[o/�,� �B�ьR�&��Ŭb<Y����g�oqq�'��N��e7o)
�r�T�F���P]��1�������)���Jy<]�g	��c_3���1��.ax�Y6n�μ��k��bDU��V�ߕҁa�����#p���i��IAT͉7%6p��2�\�u��k���uT�$��՛���W�19����Yv#�P�LPU�I���;�sE'�z=T� �ֆnQ2A$h����|���հ(*W��?��^�A��V6PIO���-�>�d��t��}��D� �H�Q�*/��R�3b�/+@H���q���?��M���>�g���K/��։=b�H-C7ǘ �޹3&x���2��*�A0[�Lfs���"���(E8IE�\�R޻�>^��g���a(#���c�,�-���]xx���L�G`,����fcK��&9:�x婪���1ˋ�!С�&�����Y������p�������r/������K����P*�P;��0Jmp�B��Y����g?V��S�V����e�} ��SR�|P��Ե�SU��;C�}wB����,��+V�l{W�w��g���#��0C���!��2��Ɍޅ��:���[�	U�0EE�JzW_B���G�������!{�C�dc�?���^P��GXI���,�S"�Pm{�8A��ŕϽNk�ƕ\Qpr<�(
�Ŝ�(���M�˂�x�E���:;;�y�||��ݏy���LO�Y[t���Z���I7�'��g�s���&�Z����i@Eq����E��qR���͵k�1���{�'ǘ�x�ͷQ. ��Zcc�&���O?bMI���7�ϿF�>W��ٟK���S����)qJ�)�e�\Vm��vd�Z{���W�cms�%j�]I��2K�stw�N���3��N*��GEk�'$BaǢ�IB��wg3����ڙB���\�qHw��n'��i��y�V^�%�]�ݡ�m����J��X��ziU��:��b� IB��:_y�/��ކ�����}��x��[|��m��{���y����FDe��j�?��k	�	l�����"P$��\����]�`��?a~�I�p�r�����?�&��ptr��������Ṹ��7s�6���AIY��(PT�m���ʗ<�}����@ˌX�1Fe�BS
Ci+�Y�6դ�M�����(<=�b���w�_�38���Lõ:{`��0����`4$��u$q��$ؖ&:A�b ���(A��5�}�7��.�����}���/���ŠZ�&Q4��)
���e�/�$	Ëp���M�pH���8�	I�����4��jj�$b�j��C����7o�}�̖q���o����9��mj4��H��S#����S� �T���g1/8><d����i����ᕦJ���|��|�����N(�֙F����Ӝ��鋈#[��4Ja*C�!��zC��L����K!���'�"$ΰ��H�k4��z�20�:�B���2�+�-�X��S�R �o9��xڷcdw�?*S!�o�	][���P��U��Q�0��t�q�WZ�]��;��z�p�L�����ٜ]�<Uqw��n6.��4~�yn�/Z2^���f��ھ�����=�7����{2Z��Ni(|�Mm�������}7_D���L�xYD�lJo�֯_��5�|���)B�]��I2�Dihu7u�v!aqu�� @�t�֮���u4�!B�&k(5����:C�>��GB���8o99:���ch��h����1��3�t��s��eq��"�%�p'���dQUTB��o��a��`L�Ϲs�C���� '7!����v.�D�3lU�Ӕ��))� �}�dȸ,�8�]Z���/�dc��~�D��+LQ���a�Mݩ���R�J��Y�i���>��8����pto�_��qF��\0o,�)�ޓ�Ȥ�E�x�T�"VU���S��O�:-y�������M�t+#���Bh�UUE��O}�.Y������2��-��t�v]�aZ��Έ���� M��,K����?��g~��;�1���bN�ؕ�"t��C	��3�2"�3�2���$��k�q�[����y�����Ӄ17��y�O���k��U��g��R���j��{�k��и���������T�RKI%<^i$ANus}�iY@ hU^ �-*|S�Ċ�6�M�oj�2�49��H��w�M�(k��z������12�8[��C�%�A�P�c,�"/��!�~����"M�%�a��l� EG c�.�Έ"�H���>��d�>��� {=\]1��br�j�#b�P,ʊ�l�����}f�����MN��,�C{ERU�霩��p���Φ�����<|�W(a[д�.4{�8}��{	FB?�a[���,⠛b�����<�^$�>��y��D���b�HQ�Ф����o<˽8�l��~�9����������d�d��-�}�9J߰��!��Ƀ]�{�l�Q�܊���(�8T�@�^	H4h�Њt}�`�������-Zv�mϤ�.�J��,d<���Њ�y� ��[l�lAhEP���(]�u߯�v�u��Ë;��j��� �?#�.L+�f'5�|����Dj�hgh$�uM:�n�;���\��L�ѻ��x�����g���Yv ܙmi�v񎦱\�7{[����G:�aS�|B$��5d�EU���CT��*"�l�
�Z��{��x����'$&N��%1�Jpb�#dL���?f��9Ν�F:���&�S67�E�8�i��>��1����XL��N&��9e�`�K���B&i*��!Q�\�پ�iYr�(���5yY��lG\��"s���#�N8||��b�M��1�|�4`q�&҆��F�$��`kff�,��[Y�G=��~�7	_;�A�ޣ:=�� �j��<�)��T�Чj�7���g�P���V�@�-,��܋78���98�,�o��
��}�σ''�����7e��l߷۔ݵ;љ.�m�f�;�C��4��$��/˲�>��!DplEp�������nĲ+н�1�^��x<&˲e�j�c�A�����=�!�d���o����]����Ǥ6�0�Q�nZb[�ujk�OI�6)�)$u�p:ͩU�/����ǌ��_|��W�MflQ��	�������p�k�:b"��h�����GC��.\�ĹKW�'�y�#��ޡܺ���"��>{{�8�{���]����c��57T^8�E�F�Q�����e[Gl�ŉ�.rR��e���: <U0�{}�j}�$�����i�-��&OȒ���o|��ܿ�}*��MCTCR;z:&���$Ɯ��w���_������D9���4��W5��ќ�H�h��,L͢��g%�t��K��O�8�,%�Q��ل���5٠���R��&�g�����H��?K@����BI|��X��,c^F�z2@����t�nJ	^z�uv^�<��YK$>�3�opp*Y�/s���P��c���ο��~�_r��>޽C�4;WoP��<:=���d"#	(��Rzd$1ґۚ��(S�xlm(gf�2�kE��@�=��]�o�93z�ƛ���=��H-�-\C��J(�3o[lC��r�-�8���2Л�A���҇@ȶ��g��*�P{PI��A���!lVD�0X��ܙv�o+��sx�|޻�w8'Zk����~i.H�_\xY�C뫼ҡ�TŖ��n��^��1��A�@i>��O�{��\�z��ׯ����`�z:%Q�����;X��L�1���Q��[z�2"�:MKCa
t\q����א����V�ސ�\����-��\�֘,����o�ҭ��v����Y��oA� �R��&�/szzʼ�Bb�!%��LJ�����d�}�D�:\Ԇ�U����M��0�/�&)�7��}����S�R�����oo���	e>CkA�m�3$��Ո���Y`�D�E�*4�7<HL#ͽ�K��o����>9���l'��RP��-)��9[:�C�FK��#�4AS�C�"�W�z������N��(Pqry�x��_�$�č[���҄/�k�<���;��dQ�]�taT
I#Q[�!�����UW��_���x֒ �n�&	�s���ϖ���pA��]B���t��e�{��.��A�jj��x*��ʱ�a��E���_��?�C�1����;w9��Q���dI�o�[ Y�#�ȡl�IT,4�$6R��{��}��֗9�Q_�Ʌ�@�'8�@|��?���U�}�s\~�s<��G���Fe��.[���op��͵���[TD��G8�37���M�EE�-��!�͈�������|̓�w�ܿ���}FR����%J8�pD�$I¢ȩMC�Ҁ�{tz�|^�H��^���/r���x�x�����,`l��}�z��Ҧ����Z�,f�>�My�.z�(�)E�g��#F2/j�lDE�h�����fB��P)f�6�/m������9�T��D3�`}}��\O�����{@�(�݌/��8瘎O1E�ɣ=�3dI�8kO�����۔�'`mA:0q
�3d�J���9Gv�2/��4�#f'��}��lG���JXo������5��ןe��ќ�풙�}�?���нsp�
O��[/]����I5?���6˸z�*�4���K�yMl��Ƈn���U�`�&���1đ �
W��((<�:��kq>A �;g:��\���C�����}���H��xf=^u�X�@o�1R%xQ"P����eɿZ�V���ګU�J����|_t�|8���}B������EK��gc��+�Ϫ��W-�)�x�=�@��m�(���/%R���?�2������a�i��"*�x2+h�&J2��8���X�XkEYW�)O�@{�M����imp�CX�"&�\|�&��=�mm0�5����Q�{��hf5��Q�5�h�~�n����y{��W�_�y��K�0"�c�	nM��4%�� :T��hĠ���� ;/����,7oG	G�'����{�T�B�J�U�C#��FԵa���ߤg�����%���_��)�ia�m����z��������,rUT�|�J����#�J������ݔۗo���=>dNʕ�_��������G�?~¸.���4DB���b���)x�ַ򻬎!V�ere}v���b���J��s��zZ���k����n����9��\㨋�Ǐ��p�c�v�!c�_��q��Z�T��U8��yCH�=^5�z)"�T�SI���o�~�H~�u^��94=���)+����n>�:�[�㋜��?|�}�&�П�wl�p���(��K0eAv���L9>�1�҆[�!u�3x0���]����}B�ܳ\��"$?�d��@1��=�s�ݞ������8�<��<�?�Fr��s�x�e�/]`:>ac�Qn�y^���8�]�a�}�7G�=f���'�XIH��#�AI�
�֊���"I�}~���)�u������x�[����������,0�0�ϩ˂�阫�;�����d�_����$I���.��~�x�K�,�$ƚ}����"l0��˜���o<���h����a��J�C�H�dI��c�VC+�ҁ��f���L��)�� U�/���7�D?*h&xp�k^�ڗ����o�&��CO����d�8�\���Am��DhF�J�]q�O�A�������B�):~ƣ*>�I�]'���(��M;V��Q�Bi��g�g�g]W�%��Ӂ���OH��r`��z��~��>��|+γz�u~p�Rз�E����`��0��bI�;{/Ձ]V�\)y*q7�r��/1g}��W��
bVh��$��^D��j�
���H�d��W6���E�8��4��M�*��$I2RS�z�n,�X����ѣ>���ڐ&�H���l����>Y�Q���)^�J@�(��4� �+Kʲ����$'$M�P��hO�wk��4����к===%ъg�^ekg��sȲlI�R2�M�T�v6�6�X�U~���K���l��y��_�l�z�f�^;ǯ���y���>aF����|�_������'�[l^��ܵ�B�%�2Q�p)O�%����0^�(�(Ix��r����y�P45�_qt|��'O�I���t���)	-v`y]��<������r]~�����2	�~9����p66����;-h�+
|w@�Cl��?��������pt�|��>�:_���xQ��kb�����/���Jy�ƤY?�]�����G���{<�l�W_"{������=���9�R%RK�W�����B5�,��i���=v����[/��=���b�`����	IU\�v���+��˷�?�s��96�]�>���{��"�qH���c,�֚��"M��3����s���x���x�)Z�\�|���y���4�6�B�`rJ��(�
��A(� 	*��3�(��ϙO�$2b��>��J�_Hd#x�{������{�P	����b��)�%M�i�g.4�����8==���akzҵJF�����Y��"j��=����sE�8s�g�>��4xoy����!w�}�\��Ō�,�\[gm��_��c�Px�C>���    IDATP1�f��HQ�|���ٹq�k�|�j�2�u��e<�կ�}p�˿�-�����G�~/+�`C��
T�[�*hx!��B��R��r���'�OG;yX��ҁ�W��?u�a���w�ݝ�����N0��ﱜ���ç��jumY���+U��˙eWi���:��3j�o��ُ.�y��S����34�<���Eh�ϵ�}�k?kn�B�,�=����̫	���~��S�e���'�5�74�2oj�8��Y��Q���%MbT���N���*��� +{��u�kk��Om�8|jӠup��OBPo� m�4�E�X�\�i۸V{�W�ֿ]x^b��M�ꪢh�<g�a/�x�q ���?5��lpdr���-��4��mm�H)K�#n����{�f��-�p);���^c���{�=n�)�k�{�s윿�}�fUi;lf[�K�g-����*YO�n#z�Q4G,�akm���1��Yߺ�W��:�?���%���f3t��F����D-�s�K���W+��d���
��� >@������/�m>��˽��X�V�����mr�mh[%PR�[��鷹�����>Z*z�b�w�)�FH��m�J�6�PU���"{C��q���������y}J��+̕།��������2ɨ�[������ۨ����L ��.��~���8�ҋ�x���׆��c-·�����\�y�����ѿGF������)��,��	n���,��k�{Ȳ, �F8H���j�6�I��(��P�9;Ww�r�"�ل�tJ����9��b�h�IG��ۚ�Ԧa:����DJ`�WX�H�}jӰ-+b������?���?��� k
�d*�+�H�kO�T�$���ܹT��z�����46Ŗ)�N�"�8���\�*멬c^8>��w�=�q�s[�/ao�l�u�y�f��ݝ���e5�l������,*�$���K���c�VTdDf=QAP����XFXVcɖ|%]�����W7�z�k��Օk)n\�sw��^s�1����$I2�kW�N�ǣ0o�g�E���#�Cn�����9�;���L}�G���r���]��ۈ�&�W���_�>}u�%Ʌ�\{�H�r�z_����x��H�%?ŵq)�Z�#/���8b�ϭ���8�"��cA	��ò��r����we����->�A��
<���<=[`�CX�V[�������c1>p���ъ���X�=��䳺9�np��)�ǟU6ѝp^v���F ��;#p�s�~ޣ�l��h,C�J�8F��Ɣ��A�`�ሬ'����qLK�+
1b3�p��)%q�"�@�45��G4�!��RX�^�e\�y�cGGGHe]QW��=٪1�jb>��k+V+8E�I�2���֜���ЪZ�`��Vt$�~׵E����.�a��4S6A�ɒ`�aJI'_Ct�x�w~�[������y�����p����W>ƍ��!�׼�W���ɯ�)����Qᮕg����只�W�I�\x�v�u�b6>��K��H�$q�Z&�1���q�+S���$崘Vy#[2�B�1�M��W-��Ž�tv[l�359h��Akq�R���{���,�je���L�T�-6�v�Qr	g.�]�ch�Q�ư-�2��X�ٻ�6����8#ڸ�����Z-Ћ:��|@c�XS�(�dK��(�s�w�u�6iz�Ym��x��<�q��)�o����{�ݾ����݌�BN|���_z����y�h�o��7#>�O�'1����6�4� Cc�4 ����1��#�1W�\'R�x
�o�W��D+���{�y�a�E��q��n߹�|2e:�䱠������L�UU2B��;�ʡ�����a�3��qi����0�9q��s����^c��mTQ����~�����=ύ�W�E/L�XO1�RNf̧AQJ�����$�8"%���.�L-HK|������ӢjUP��S�&83����~�*��-�7��������ݷ��__�!��IW �W�'���|")���k�~�:4���~�c����ظ�,�'�����߼̅�ߡ:z�����p]up҄8���DYڀ�SU����4������zz~V��������=��}L�U�����I�����}(ϟ
��� ����g�Y:��^�T���p����[���nI�;�}xS�s����W �E��l^_�j)ֻ'Їż~���@Z<oi��n�e=A*�j$���#4L��� g-6��H��#r��R#�[1�Lp�����XS�IE*=��[ϑ~SяD�����=�'Ǥ�g�V��F�$�ڀ�8g0�&�F���{��M��ČX|5"\+��L���$qK�JӠ}�|�Vx"fݥ���՗��� ��pg��	�o�BS�q�Cz�&��e�����&�~��?v��?�:�ќ�ل�|Dck�i2CK�m������Յw�shӜ�{�,�����bo��k�NA�L�f��fF��26�>�PUزZ��'*��A��_Mb�_@«��T
θ���E��k\$�lPcl�)1�i+�3��"�^�.��g���N9�<����������9�[Aˡ8a#�Ȳ!�:�VRI�����hD�E��6���^�z+��4k6/n��7^�������Y�t��^�1����[�����Ɍ��S�cd��XNw3��˔I��;ֲ�{?}���~@��ܾ��n� K;�M�l6a��#�|�M�ׯqtp�������{c��5�b6"^��Z�wz��c�dYΨ-��	J��K]�r6e2Q�%���&K&̋����R`kA?�$B`�
W74Uh��y����(Xg2F�`M����e�qݸ�x\�FB��{������Yo@�$�I�d2a6+���FK��!Qx�`��K��0���|D?K��4"�y�^
l�PWk�xZ0�k�u���dFYΘ�s� �=W�\��������M�����n���YV$UMBD�R�)�`����iH͌ٿ~��B�*��v�ؗ��J��|>��?�w2�x���`�=_G	Q,i���*�J'�XG��P5M���$?�������+�E�^����<d�3�} �+��{��o��hQ��O��
��U�������xRa��8�B�,�Y���LPdqb�!E � �'�~�Moyۖ�b: X����X��*�?��p@)d�Z�g_{d)����i��A��H��ł�ݔX
�$��(��0��!�$:K�\��	�	��x:�9���/�� �"�>�R�%�ٌ�j�t:D*�J�3���g��u]�Ҩ��P�g���uSA�TkI�D4�n]�i2��KW&�2�W
>TE���ˤ#H�:��$�b::"S�^��"��/�2�����A�5�U6�]����wx@)���D�FIO탳�D�����|�;|�&�U�U�9�(NjE�t�׎y$Ȯ^At�D�ьZ9�j�>�W�"��.��\A
D�E���WoV��'��k7�+����童��ς���r�����@#y�s�4����錍��+&4�#�(��di��P�mhR`0�� �"�(���jt����3<a:+�G�s>x4�4%��!��#�O<��;�p�������'�� }�����2-UɃ��r�n��k���XY��qA�*f���̽�鵎��鈦�H���1�iA��D68C^�x���[H�[~F5�q��6���l���X__'"�����ho���c<x@�X�(Fk8>:m���p6p+��Q��뚐�;O�$�1�VN6 v���}N���&$Qޣ������XRzC	VB9�9i�wH�~�O�4����t�bG1�NB{'�i��:F� v���c�ݰ�!	5��%����+B ��4u�p:��(�<�V1Ͱ�<@צ���+�<~<��׆��}�����sz8�����1�0d�9�����+_�m�z�X=�#^����7�>x���.�)�"H�Xoi��M��5Qۧ�&�)D�o�u�g��*w����]�!L�%�Ok^�()Ck���vΡ��b3Y��<cpK���������Kx=\�v�#��yZr�����^�p�z�ߗ�y�:Vu�/b��Gۦ
��Hdx#��7-��w��`���PA�S)4�������8dG��֧��IK=���E�8F�/"�8#�L�
�l\�$��j�r�X
d�!K;zkˊ��*�4���0�����8g����
!Œ<*߅a��
�w��,���A`���Z�eEQ�4y��d�1�<T�n�A��xWUx�ё��&��Svw���3�3�����2��3�����O�S>��_���ӽ����GDN��!�s+B@+D�_�|����W��y��h	Vh��"�v�O�������q�{�}����=��)���Ԝ	�<M�y�/��'`�E@^���Id�B;�L�E����~�Z<�i�gq�3Z�<��.����3*7"N���@�a֠��Ne&�����΂:�d���"���v"|]0+J�|�<N~N��N�q��'�~�^��wH6���a{����p[����C��$��!��b��M6_�$n���d�\8���9Y3�xx�h2���P9�m(��C�՘��7(j����6���ϐ�1�dƟ�ٟ�����~��x��w���~�/��o����QU	�+��#��U�x6G��H�^��dƤ�H"E���u"��G�$��L)�C��4��G�$x�U�u-Cu9o�:T�x��):���{8�#�{����yO�3 V1�+��4���	�q����Dy Ӗ�5i���L#�& ]�ې90ΡZ�1�8\e����
���,av2��p̝;w��1ãcb�k}�(�����xF��8g'����f���(镂8N�6w0ij��x���&g�<t���fVp���+Flݹ���YB��4&$�M���qΜ�N����J�?�<MY��},{�+�ku�Q���r�+�w�%��%��_YV�pO��چɦ�P��.��;».�Rjh!х�N���O�Ow-4,�i��hZ��`-�{ჷ���}�Bx�=�P�/�o�儍y�I�ZN"Bڶ
X���â�L������n�!:�~/}�
G] �����PGJ<7�e i
qTR�"��f���O�ωT����TA:�8�Ɇs���?�3u�X��$1���>Qa]�|2iq�2�4��{��l�d:A�NF"��j��38[��z�S�`����Ea�C�����ե�)a<�T�X�9Hc�t����k��`\�4���~�/�}���y�������&������l�X:�����$a��L\� ���V㼠�6D�s�I���"(*��� �9<���FR¤BuR�tUʤ�Y�q��7����w��Y��]���@��9�L�5u3��B�ɺ�1k<cY%
U;0�ZA�D�UEACb%���ƌf�Dc�%�cb��`=�0��fadIj�H���k�nƤ��eT�̥8i���j�)6�N@|I�=Ro�V5�VC��5f�2�z�sc1&�.J<%R��Gb�g���5�@�$��K(f��ԑ����uCS[d!�Aق5�����h�ᠮH�.׳��	�bF�3�;����sqv��(��a\�l����[ě�<���M������&�������v���TUEY��֐T�(�2lP�K�8��~��>�⧨��p��g��O|�y���^���%F����߂Y�BДe��4F����He�7	�K�G�����*�i�2��4'S��LEC�A�j\�q�
��hQR�v1Z���dJ������O�����̊�r� �%�ِ4YH���51 M2F~�kD ޵{�u�"{ 8kq
�	mY/Hb�@T�?9�(+.\�`�B�$�A@I+�7$��(�)�!I�뒵<g��m"7g]A�OP�a���D،f���9��	�74v�H�Lb�-a]tq��8������E+E=�����Ѹ�L�$&��V������<���A�@*��J�6H�T�V��F�[�<N�b7&�aqm��/��PjbJ����"�AF)�*@�K(s�-+���Y�p��������t�ھ�#\� Z�!�f�o!�%�B������c�7�Jx8�--��'��G����;ψB �BX��vW���i�F�"�+Ic�.C�.*�hS��	�q��u鶴�8���G&	'�[iʥ�Ϣ�{hQzOB�zg�,�g� �zrrĽ{�8�Q%��%4y��jHK7��Z�@��&�S[�u5�L�u��P�51r9C����6�=�<qd���{�1T�W9ts\Ull_a��}��;����?��\�elЧ���p<��ʷ������?�PL�fc6�M0G��r�@o���ԧ�����>�^�\�H�us\��M���I|JZZ��'�y��?s�=��c"�b�K�.]d4RNf���t6EGq��jPļ1v��.qR��:��0)J\���#cEa*BP��8��qB!�Ή�.�M�#-��ݐ�&I��,�2.k���N�a6�s��e&�o+"Q��cr,r:G�"K��L�'��$�����	��k�r�*],��� ��0�$IЍģ�Ts�'3杘��dY
Y�� UF�G��3����ݜw~�]����S��C��p��}r�o_���̚��h:i�(�z����T5���O��I������kW��/�R�f�ol #�w��9<>��>�ljPAut:�1X_�����h�h<�i<�>�"�[̊���y���	Y���3M�d5�i1��5L���1qq-��gi�����`|TǔX$�e9����QM�v
Ӫ1.���V�iJ]m���1���Hb�M��%�ښi�4 ߮QOCYW�ʂy�<B
�sԍiG�$q�`]�6��!5ND���C�y�n4����C��E�)�1����L�����x��y�MT=��� o���*P&Q�,>X�j�Uv%�'\�qgqpu�Ї?�L~2>�����d�m�����X���kG!��)B�{�%�~�9ƷB#,���p���X8�<�'xr.7�Ǔl�6̷�Y���Pއk��)�&�����u�]�}&������{2(,��L�=S��������Tٌ�w�7��>�pDQΰUEGH�1��*�h2eR4�G
��X�W�n���ú�)�y���X%l��I�>����z=�,C�*�vy�t��ѷI��0��i�Q�lt;\������	D�#�����HR[A]�E�t^��*�-z#l
BIDݠ�0O��}	����Eتfv:�Ae��R&U��x�����潝ׂ����.P�\�f��Ox�����c6���;?a3�p�0�J*R�����xHx��Z�W�1joi��+��Ԧ	�5Vh��w8b'Cg)W/��w#N�?$q��.����o���}��w�Ҍ�������g��98ݣ8>ft�\�*�����&'e���+|���j����샇H�f���8i���h�Go���T�D�z9�I9ј
kn�z�KWo�{����]F�{�Y�t{�/|�78������0:��Mt}�Ƣk���L�4�+�i�)j�����>�/np�p�Y�@h�ܜ���iIi+�<E����2̄��c��>qe�;]�/^d�a:i�����\}�<��_�׉�5�KۨT3+�4�&�?��:j��U��w�[���J�E1^{�ց,�""!���������:Y�RU%�{���/q��M~��Ox�����{4�0Mpx������_����?���9o��3^z�_B�e����rIZ�Z��9
����i�x2��%=���19>f63hl�w���.���@ck��N8�
���GH��K�w�d��!��@�5!�Ǳ�Yɼ�Q�t��HF͛�"��=v��/�YQ�x/"��[,ec��#�1Y�rR����D&��;'p�bm(��7i�G֋��4�s<EE]��#��j�͔�ŌA���#��υ_�*7_�����K_������b�V�$�QBP����g�`�ɐY    IDATy��)BPv���K'��ں(e?Z������fO+I��o�t�0����WY�E��� ��jo;��W?�\�"V_����� �'�����'9���b�p	��6�A���g_���W5�=gH��9.Lo�}��քˌK�8A8|&)WE��N+�A�����&�防,>�8M�ZGa(E��DI�:��B�\C��AJMfDY�k7ﰶ���������fvcC?�ʍ-����b��E���qzt�����#J���ÂC����y:��J�ӒyY"�^7�)C�X���:=�e4�Q��`0 ,����f�ڔ�$� ���5"�X�0�<ż&�
gj�ܐǚzR2�xm�GG���=��]��o`�ǫ�Q2EXl֟Ϩ?��2s��~�k�d��y2!1�!�)H#*%����|�+>��pwDå����{Lw�q\�ڗy��B0����o2�?������?�����ɐW^�g��2��'d�����lݺ�����k��ʫt|᳟���N�d���!��.l���_��H-x��AO�=x�K��y�4?/�	N��:�k��;|���������>{��`8�7�7����̬�����������˷o3��:��Gd������We+.Lt"��Z������}J�=	���l��k�����|�k��+c}�Fg�O��A�`>�yO5���}���M��}FUæ�3ҤK�R�"Im�l�K\dKe$Y��`kk�n��p8����p�Ԋ^'��Rt���s�Xs��%^}�u���#�QS�e]�PH����A'�S��4�=�?��rz2���(�	{��A>ϐ:$@J�IYU�u
ΗAz�B�0���l`�/R�f1�JS0�M�F��v�b,8y�'������,I��ӥ�A@��7�:'R�i��@�J�
�@�WZx���xEP@��
���lhM��BOB�lp�K�,��Q:B�	*IёFi�L5&Jȯ���W�+��)�TD1�ӄ��,�()�]�"Y��r��w)?���M9�-���@*�.$�m��˶�ݪ:.{�"����-�S��'��2>�r��G�R��u������Xk�mt|���be��-���Ӳ%��<d�$�H� ؉V�WĊ
�_fyjy#,��a�Rg������V'HI:g�7�9�Q/R��[eҷ���Z<�������_�{�����t~�w��ȷ郀Ѩd<}���y�N����8(�!b�H�,x�ԁ�([�K�9!J4�ٔDK^��g���MP�ئ��U�q��^ଧ�*|���)�NJ��\��b������A'@�Jd��d��V]�d�s�u�^�ù�������hX�� �b��xa��&02��I2X��X�d��˒����3�cvd̍/|��������������p%�Ƽ�?�_������������_�w&�Sd�I��L]#d�
%�2~��[Emg����D;v'�hG#����i��	#Ar�&W��o]'�-÷�޷��t��Z�ǣ��Ï��%��NY�sRc���������x6g罷�{��`�b>�ݟ�ɻ����蛆���r�?�9?��OP��PL����S߾F1�Q{�l:a~z�h�!ۛ=FGCNO������;�X��F�	�k�u�sF;�Y�t�B�u{\��d��ؼt���|��ь���q}k������v�AD`!�d��c�Ǉ��E�?S^����J��Y��2�U5�;��.���O|:G�P�55i,�e���h��Y:Y��`���X�K�i��t����:�m,W�ֹ�}�+�����I�$������!���E�t����@,��������;�i��z�ݽ�@��:H9Bˈ��C|�Hy�8���-I�ι�{<��z��n�}�'DZR��7�ASZ)A���q@�i�[���H�$���'
�e}P����:Ut��M��8Ak��} �1TՄ8�p��Ҹ��O֒�-�ϳ1셔�s���8�E�-��$d����L����BA�wTKdUaM*�l1H)q�;��m���9��^$� 1�'�czL�����c����S���d���HӔ��1ƅi'�[�|��]����":?!F%]���q�oO�?��0�$��]z�Jo�c�A[���.g�R�b�Ћ�� ��:�ً��������旿�-�p�XlqX�C��-�]D�@;�Y���	�o-e3�!�^�
[R�<O��^������O[�;@��Cz�������I�i,˚�6�ź�f�׭iۗ3�F(�!��O�!�47o]g��6�8���HQ�F�+$�zʺa8������c��!n4�99����y��y�p<r�R��\BPVQXP##qR�v�"~c��448&�`�p��]���#jk�4�`o:<=����g��I�%�"�X����Q�F�s�ӟ���l]{���<���N�Q{���^���˷��y�HF���c���G; �^S���V=�m���w{�^p/����R���(�o��;"��!���M�o�Kvy�T%tֺ��a�oP�'Y2/��?�����?O)6ӈ��c����
S��V]��(�o��Uv�S�pm�#ʂ�4a��}�����h"͝�=����Ç��/��!�6�sz�f�ۥ��H�b^�o^ANO��1��姯�ʑ3ܽ���لr6B65��:G�a|z�����g��D��C!�Wq9�`8$jR�(�p���cSЌ�Dq�*�l��	UQ8oH�jkqRQ�Ox����s��:S��ҟ�F��N��D�o�/�_��?&_�c�E�P�q�b*���l]���z�z^�u�
�����92pgYU�����<õ[7���孷ޢ��D���DR1��/����2N����ܹu�+�.��^x�,�y�x��a�F�x��@Ɉ,��usz�^�6o���a\ʹc�M��x��a4��0~k]4H�(����b�,#�c�8&V^)��ԭ@X�� ;�o�gIKR�ަ��N�.���7A/CG�ZG�͇Ϗ?{��"\�
�uMS/}:��кQJ�Ě,3�X���X�XSl[��H��B�PޑV_z�#�����f�gos�wo�IKÈK��e:�ܤR��@9���B��`N�D`֟����^����Xa�Z��)��j�X��͊v�Y��d�i{�Xr��H�ǹ@�xC/Crz�����lW��rg�܇����� �s}}Z�\;B C���`�[>,t8��ϯ�ɶS �b>�`��z�O��T���ZѾ�j�·Ν�x��w#3�Bā�В7�C!�وDX`UP)��r6����|�v%[���h�6�أL���ɔyQ0�L�'c�����S����<<b��!�x�7�x"�jy]�P�$Bjڱ{J$*��z=�N��	dg�ƭ�lnlb��(]�������`:s����t�L
E1�0��!�	�J�>��F�Wh�|�9�=s������7����c�}����)w�O��<��D�������껯a��Z�xA���8/���GT�އ1�����wX+� �<%iK�{d3��������D%+��`n*R�I+C���.%]�f�T��<l�u��+�s��'��^�q8��G�r��-�?�d� ��(8-<���<��K'�g����%���-
�1��F{ŕ+W�r�r�1|�.�[����{�GLf�?�܋$�bc���o��ostz�7��;q��?�����N(�C�|��ko���	Jg�6A1RI⤃B0�eX�ί��Z�8�B"Lh�Ԯ!�$҄�ix����c��e���8�TUMGF��ϼ�%�[�w��v�!��;��/x�]D��r��-6��)�MiIR	H�
	ݼ�p8��a���l�B��w�ec�2Y֡��t����)o��U>��}�R\�t���S�vvQJ��v��89bMIw��e��7�7ll��kʹ	
��C$0��D�
X��H���^Ij���-#��A�/��jH#E�g��ֈӈ+�/���I��xo)����NN�"L�"�!ip�XG�ч[d��T(�8�W��Z�KE��l]��t������hL]�qR�e)�,02��[Cvl�P���Z35�x�ݿ'.�w��oy�ګЙ��;�e7�˕_�5>v�*����"���eY�TfI�S^�{�"F���������_��}.����d�޾[�Wci������o�R�/Z��^���?>=�-z�*\O�罷qV1?��_8z� d|x�M�d��>:!����g�^,�����8�!�	��+?��%�	��/�z1P,��U�_�Th�F޷*Fm�7\�t��t�AE�$���	��Z���E���u�j^RMG�R0�����;��%�9�8e<:����x���q�A� ZӸ����'�MYKb�d�('�A-$�����B@Z�_��@���q�x�]��F=�U�I���>��8NpR�]z]�3�U���6es���q]R��4e���c�O)DE?�3zݜf���[/��/�e5���gs6���ɔw���_��?��/�n�3?��K�R���K���K�G 5��ɶ���_�9��FX,��N�&9ESc��n�G�Ԥ�F�F����n֓jOmas��d4����̌!J�a�h|J�e0*+jW�uB):q��e�$��`i�[�<���ŝ�êF[C'�L�Zg��p����m�M�/_�2�X4�+�[��Ir�RuIk�������6�)����7��1u&I�WWx�Џ4q'BH^��$a�ux-�w�j~���G:'�<��KT��EЍR��~ i�n��ڵ-���xg�3��5��:~s�Bϲ�*WЈ�5�a�&'c6ok�<��/�$�,ToJ�U������	uYᜣ��2X�39>�������� �v����p�!����_���}��p����?xĴ�18�V����1�5E���3���DF� �P���$y��e8��"��8�X�-!��uMYT��s��_;�r�b]�:���}�67x�S����=r���d8���{\�z��4�q�����C��.ei����R���Qu�S$$q�TxϠ���ŋ\�~��~�zgʚz>c>nh�@�(��ABYkM����kE���o��^����X��w�D�aT��.�sìz����9�ے�ӍJ'�eCY׸Ɔ��)$���ʦ�g$9%�-(�S�����DP�[�G�R�ZX�/��I���;�q!�S_s��ڧ��w)ĘhQ�Me!N�ib7��y8jZᕂ��o��[V��f	_�Yx�{`
B�,�B��A��혝]n�
%"j���	�k^��@�S�# |�W.�ʅ;�w�J>���ZO$C��hP�M�Ռ
I���ɉ�`M�H�Q��w+�e�"<s�01e�K�
bs�i�7���w��A9�h���Y|A�ykZ�-����U�#�p�F�Z�amh�ԍ�J��#���Fa�7�(Q������1[f��W>OOy���lL���n�10%������G{�J�sME�2Qk�8�'̊#��|)倆*3D��Q�t*��>�E�є�����R(��$��0�'$F���l|�'�A�!�"�ʒ��6w�}�aQ0{秘��j�n�9��"�.>�L�[�2��5t$�����d)�����tdM��N�Q�TJ\7P:����է��ȣn^�����#6bn�\�WΘr���S̏�f�V$��t���R���(�y����%K];��w���$�Q��4G��hNy�IlMY��)Ӄ�̇c̅u�$���w�1L�1:� \��k��WX��6���bP+$%/[R#+���Xop��xEn$����߽�s_�
ϼ�YW�pZ��mv�!?�ýW�䗿�En����o���>ɘ�zC�ݍh�l#�ڍ�k�f�C(�1-�|����1�P�&$J����������v3��X��%[6��t:�VB��rD=�yú��L�Z��k@Ť�.�>s��{0�N�.�hN+zk��4��M5����f\X���0J����V%2r�DU�x�H��N���KRƲ��,�h�ڥ��N���ŭ[7H:9�9�q����T'�Mح�S�ǀ;ƛ	J���d;�Q�0ƙjE"5�k�KG�H��cTW􁍵ֲ.�l��W/q����HΧ����h�w�c�Jht��6$T$1Ra�+k�͌:�tO*�f�ދ�"]�fm�ar��<x�.����2��e>�����r�WN�xD���UBmTK�8a���h��P^ Z¢}lE@��jj�l9X� �Hv�8��İ"'�-�Z�� �2Z-�-��@���
�[�P$����|(a0*	\ν�����4W��O#�����p���V��PG����gF�#%���'����g-$�J�!x�y�U�?'K��؏�y�!��)&�R�	�xgt�b���U\�2,Z�i���8{�ɲ���s��Œke���lvSM6M��DQ��F�@�_l��"
0�7���� c�`[$����	Q#����a7����=c����pndfU7i�HDVTDdč{�o�.2�UC[�8���C(���<�*�m�RIs��M �!��px�;�F	A�|��-18T�tmHf��!JB��g��h�p�y��s���{�g�8�[�R�{�LZ�JQ�E�ֶ׷ϓُk�h���f������r� -�p,��]�˯~���ʽ��6�S�⡵t"b���䙧 ӔM�Y��B`��Nn �p��x�:}|�d�Qo-(�f�(�6�`{c�����Ss�Z>%x�y'ƈ��@*��4�c��锕�y�G<z�M����ۣ�a)���.:�&6��>Ǉ�ƯPJbT��dJ�k��M����6���טh��h�ɽ}���ݹ�W>�y�w�����3�Q"ZO��X�[|0,G���dd2�_�X[]K�J��q��X�Z ��a�iM���$ѻ��זP�!�B*��X��Ny����O|���)��ښ��K�W��W��}��<�ɗ��(�:�b�ߡ�O0t�UM]�x��ʠ��lT��,\�4)$�dP�de���	��}��ns�8e4S/W������t���4Y,KE={��0HG��HFnal�z��&���[tmM5�(v7i�<|$��j6�6��SFf���,w��0��p!���h
iP��o;�stV G���&eQ�R!����(�y��g�{慄;0
;�2麓/":�r��y~��Ⱦ�=����?>!,JS����E�*�$�e
2m0yN,3(3ΜA`���a�z�ܞЊ��dN��#N=L� e�Ѵ5R�2��la�F�8y��Z�a����W-��"UE}s�O����_���s����9����v�l�p����ԧYNr�\�8�st�κ;��.�'����z��p������?gu�*_�W�����ֿG?�N���˓�~��m��/���@�[��q	�u�!��:���J�Q��3^�K��@wn��EZD"
|��5]A$ ��R�O�����mr����Hx��O�1}��\ 6�HHu��T�4�L .}~qNi�YAn{F���Qs}�&������t�vUS�]��7�dYA㓤���O���,��mm~�Sp-����(�e��cE���cc�
���5�|�ζ䃜n�4�G�鄍��%��L�y��k{;EE��t͊�Zn��v\���k{F:C��b��Ǟ���{��>�ك��]O�ߍ���_��/}ڎ�7ߦ>>%� �I׺���^�\L�&�B.�$v���w���1���R��u*3(�Q1`۔�ERź�H@�ȏ��x��4�ӷ��+�Qh�s-�I�	�Lj�����B���>|��kr�(�9;r��;���Z*����fT"�݃���W�?x���ş"e`����������QB���uqr@�7�#oV�*Sk�\W���{h"D�6n;�'�(�D���原D�Ͽ�R������#�G���/r�Oq��������7�/�³_�/��W	F�(	�c~�7����;��|=��i4&���5z6'����ENbt��`]�rvt���!g�Gd}ϧn\�l��Ç�x��6�＃YP_��    IDAT�*�_5�~�Ggf�X�L%��#JA/s5�d;7�޺�ͫ{D�x���Y��P�v��R�z�!��)�������_��^��f��g�z������eL�5�He��D@^��`�����= fuG�i��VH"�Ct-G�����wɭ%,��}�~�:��Ry��Fr]��Ǩ<#� �@�D��Z"uN09Ս=@�]�eAČC1;ǁ�U�@2�(��h� G���ʐ�<Ԏ����>���*�x��׾������E�<�'�x�o��K_�֗�*����o�C=��/��."�h���S�1��1���t���s��sz�Gş���C""O�/b�G{crl����וO|�\��/��'����x��5��|�MD�dh#�� �8��Z���O� ��cn�"|�	��lH}��Ǔ��(p���E�0\�+?�
�v�z�s�������=��t�ଠ��\ �=�>�+<����bD��k��C�x�R"�]C��p��m{����ı�]אI����S��Ɵqz�>�(��m^���d��/Qw��L�ѓ�("M��:���cr'� )@ֿL����h��)��*/�����'k;���Tx�Q��I���o�M��o��ۿ�˿�+<���| �[=N�`R ���������a���P�!F�� .l�'��?4'
���P>��p1�H�J��չ�0Il��1��
��Qנ;~��5���C)ä�X)��ǟ�pCWHk�F������G����5��@gɍ'_���s6ێ��Ѯ�("��s��гٷ���~�o�O�>��vE�ϖ#�2��9Fb6Gd�lwFW�@����p�q�X&Бs �V���L%	ϵ��ڛ"x?8�u�?<����Mlے��%��)��$�ܢ�����gW*��?%/|�K�q�����=~�����9���d*�2�j���4t�w����&����r͢^��?������3�A8��L�4ǧ�ݿ���Lۚж�۔@XO�u�c�M���H4yH�e1��ߵ����?�{�mT^н�6�K��$���G�8{�]N��i���ﾈ���ߡ;�'���:0�+L0v*S#Dp}���)��}�==�oP���yJ����R|D:�[���������.��G�ݒ�{򲠩�Xv�m\Lj�A�*X	�
��9�傅�~I??F���Snl�O&�c��j��)��\A�6�񴀾%����('9!���U��,��4rmr����'����L�=��f��,����>���m&Ͽʕ�=�8~���=�>���p�������CR )����!�]gJ�K�����}�z��F�]��A>u�ŇD�\_����Ÿno_�� ^��?�T��,~0�C�C�4h_<R���rkQa��־IٕLٿdm���B��)�KAZ�T�?ǟ<�������]NxR?�D%�c�/$~׏�B$żH�h_:���
��d�B���y!P�z۠��T3.�]�::>���v��2�d������9DL���h�P9B8%hE`e;�q��h��Q�<9v���dt��@���u�@��l�����:g�FA�Y�t���4������̌	��|�d��lu�O���M<���'^��+�GĂI1%3��w<��w����}�ED�!�f*��@��ć�a���A=,Rb�A��0RPH���
!�u�z4� �Ԯ$yb>1e��I��k:��hcP�C�5&t��&1`��"�ئ!��9�����d'L�@���mZr���k�;�<Cf96B��s=A@�5�mX��0�eN�:�f	]��:�3��d�"�o��Dk���'��"z�h4v�'$bHd/U!���ǐ�q=�K�W�p.nD�1՘�dd&�N2M��|�Z6��S���?���������XAd��j8b�d$�G�;�r�����Yu-Z)��$]�µZ
��n��,3rm�j����A�@G��[�T(���~��:]+��b\tg�<�����>%�Om>�26<|�5L.����C�r�	���NJ*!	��x:\���+�B�������� ��(��������w���_��O}�1eq2'oz�b���z����]��;,o����JXt�&�Z�a	h�q�Z%e?!1F��,=�]�����C|�2�v������LʓHAg=�x¡J�A��"ט�q���CKP(F��"Nx�qI�8��ߧ{�>�L4y�d�
�*��@��� ��E��uu
�C9�:Lc�����Cփ'!���D�XS�׉����#�v��5RL���N��]
�5:8��,u.=�r{�2�u@�DE
1�c���n"�N�c�$E$YZ�s�K�>���`����\:9i�'�*�� "ka�8(%CX��������u񹆳��s��ɧ]��	qYg�Ck��>&B�;A4
��h~�]��S��[ϲu�:~�K#>X�zE�X!�b<!�%�Z���$J��v=�b�v�b��n{�f�r�+�I��$����'��]��Wn=K[$�������G�2hS �'v#��X0�$Eቢù+�U��JzH|i)���{������-�1�Sch�#�������d�bWG�V"�E���TdԷ\��h������,h��@���]QZ�R"�h�8��{�A)�L�c��ɾU�D�@�Q����?��Kɲ�Q�4��Q��B�^�2`��ipD"W8�*�|GO I�IפΗ�()�C�X�4�ـj� ��� G���<}�h)PHb�ڣt����B�D�B0-�D�:42͛�P�D�>�/�IP��+dJ�<�2=��.�/���ؐ��Ħ%W�����'���KE�`vx��j�?x�U�@iX�m��0��l}�%&g�j��KoF�E�:�"d%M�$e�Pdt��pNq�:�c:�:4B� �z��d��(G�I��,]MD^Z�"�I�+i	�=.��=-8����e�BQ��4��lEC��Py՘f���aNf���Ŷf٘�)�	j�Cv�G��J(���q�ݷ�����C�~E5�y�?��c���^ac����z�����5���I&��ؼ �� "+�b�-�1��*FMO��+���8���2��d�P�g�[�2���P�o���Ţ���E��is�G��3�<��Oqg�M��c²�W�PIp����]F����
�/Ų��'ʶHĐ�K]�p>c�)�\w�/`�ѭ_�����p��-<�G���'.�1x�����=�����3Z��/��b�n.��/������D���b�M1�	&/(�JA�y��W/�]�o��M�.�!8b�1�=$ܻD"��^]zO�ӝ~֢k��ŉX�|ئ���/|��C�!��X�������c
��@�1ȮֶG�r��d;�����K��1/�FWp�%D����IT�2G��)\�� s�%zK'$������ۖ\�MKa�#_E��n��=��2z"�޹�
�Ԇ<+1EN��QdFQd���Q�fւz���'���P��c(L���`l#Z�5�lo��������W1�M����32���Z�	������sZ>���$�u���>t �]��kC
���S�*I@]�I�X%?� Y����G��HЃ]l���%�D�#L�'��x/@e��"et.,e5����:��������;���w	<�iE��H��6��U�%�L�w��F�ƈ�h�qJ��q.Q1 P�A�ࢢ��El�\��>�K���Fbr
!������!��r�㯲s�y�ʜ��S�;W���s��|��~��/�;��^�}��Rh���*_��xx�6�޻�����c6�v1��x��p<?÷=J$�!��k�����@�+�U�s=&F�j����)Rkl�.x��&7�#66���%�k�"�9.�EF��lE���&�Y�M����8�P�neY������Bj�� 6�"66麖f6����L��(QK�)�������m�FYu��{�NГ1��m�?�ؚ���q�!�h�VW�eյ��f��
#]� g�]���G�с�)�\fٕ]��m<�&l�\���!\����,K���A���}R������2�����Ӛ�%(5����#(&��xg�����<��Q���vd��ݺ�̑M2�$)�T-�3B��tRA����(À�\����;Lp��1k��k^�A��x9�Tg������� �Ɔ[��}�&(�GgOާ��0�^��E=�6�&�\����3�Wn"���|D�	�a�B��������>��#���]���#Ȉ
�F8)�J_�Ϟ����I�e`��5�S�s�].�\��=J�h�c�a��%,�Zx��d
1�&��{�ƪD^�F�s�|�é�:#�D-�H�@v=�FFFH��D��1��E�#���4MoɄD�M�w��SV]��F�e��2�%�(���C;�P���
b�8zt��m"Iٯ�GdF���W�L��D����S\�L�ڀ�{b�������}���:�
Ĵ�|�e�EOӁ���[\�̋�~��dA��3������{��=�֠��I�R�J�,�z<1V�O�.�ԉ��[���Ja�����D_g�dI���L��I���'4qu]�L(t�pxbJJ*S��%���֢����%��N�R� �G����)���2��R��	���Z�)�!U�@�-Ӫ`%#*Z\�@�D`yvJe"&�IV$6A�JP
�Q�l�Ud�h�H�tށ�ĵt�ci}]>�SZ��o�9@�I����۷�>��/�*~T�|�5�`�y��*n|�kl�W�m���?����\�ԧ�u���p������'G�F%��F��Y6<#|�U�|���USspz���n��Η�9Z[s�8&�~qƩ���tdJS�'�7���g?C��$t-�pL�};��aS��"gu�@
��n]Ag
*����6� Qj�b�
�vlW#\5b���G�:�a��e �̰J�o��/�]��"ֶeF״�:�`������͛���5�Q�Hh�5�Gf~�bF3[�sM�k�_bf'���k���'.Z�0�׹��ϱ���p�T#�֑وo�n�x'�Dd�96�ф��)F#�e�F��C*
�]�mP�C���J��r��[<x�v����o�w4���K��&�6���C�n<���6w��{���ߒW�>~}&��0B�<��n�:h�+�������*[���햏�����@�E1}��g���.��ABtĐ�4���c�{`�L.�-�w�r2��$Aj�w��^�4W�z���#f�����|Mh��O�h�(KDQww�|��[D�P~�Bp��?�=|}x�̵8)�At�UX'p}��"�|D*�fFq-r�>1j��F�n��5(0F�� � O�M�d�X��L	�r�A���4���f5��ӧf�D���d^1ζ8n3�~᫼�o�[��0���c)`k�l��@�HV7�lG78�eEZ��`��{�2H���˚�np�MA���?�1��~�`�*q}�jl���<�k���L:��5O&ϙTc�4	��$�a��f6 �י�W\/�9�~R���Ɍ`kZ�=����9��ߤ���Ͽʗ��K9_��ſ�������+���ɷ7Ț������O~���w�3ݻ���c�lOir��j���p�����y	���#�1B'ڧ�=�af'.Z�1F��=ZhD\�\���(���Y���3�LS�,.sH���� F)D�J�Z��wD��OGR�\���FK�	D��W��y��R*B��8�r� F���%*HbP��-k��G�|�BK�,��Q}K5�2����1�S��nW�H��85�U��LT
�K�j�O��G�P�2�w(a�Ra���p���w�������L7hC$�3�_���oxtg�=�����g�g�Wh�V3�B#7�,W+��S�AVT.���E�����[�8�8U
��m{�M 6���������8?�佟��{��P�X��s|�d�|rb���n��H��Z�mK)V�f��3)��fm�`F
U/������a��~��ܜ��]d�{��%�ј؏(��u+�ﰲcak�[{d��"���m11�j��NF�Ō��{8-بv�t/�
r����?�<��'��G����B��l899c~|�.JF�{�DleE�1I	�(��آ���8��;��!�e�&-jF�当'{;�ÿ���!�w��W>æ�N�'zA�-�fxD�޻|�/������J�g���akr�P��}Q*0����C�߲"���"��� �мL�E���=6�\$���0Q18�(���1X�\'���B��0: �(ː�Cr)���a��<�'�z�[�y�� 2O�������H�{v�V�a
�愽O��/�ȉ�X���[os8�QPd%=Ѷ��$���bkw�W���1aT�LL��S�2)*^��K��5�o����ȦL��&ϰ�Ya�>UmB�{���ϡ�'>����;O�vL�v��rr�Ok[r����C�AP/��G�<9:7��|�+��(
BZr����}�)�]�`�l�-��h3 K�eJE�6e�>�M��G[�s��� =ݨ�L�p�:�|�dk�c���o�5Z)v�\�����2��-!�Ҍ���kP�#:G'=�����ą�'�
c����FT9;��.X6�{�/}�w��7(�b���_|�lY㿳�g?�/��o�h͝7~����ܽ��+�0��g���{�G��'�
$AE���ϳ��O��ĵp9+�yY���P��Li�Z�C�u�p�ne�"Z+r���@#�d�@c1��@�q��(�u҉	��L�Yr��DBL�����^�t��׸'v��� Mߑˤv�q�jJ)79�/��u��FI��ۭ	&���u���5& I��n�P��qm�?�/�#?�q"�`4��&�F���h�q��[�w�*����]���d�ʷ̏g��mrg䣂��n�Dd1o	Α�{�}r.��'e�6�4m��_.��O��!��>�XI
��h����{{r�yk���,�m�4
!#�Pt�eٶl��`�B��b2��ƈ�Ye�l�U�U�"SHͪ[Q�%yא�<�R�6$a��5'����������a$��DY��mKY�3ژr�[|�,�}�&��e�RD���t-E5�mhړb��⤓��t�,/��cm�����[����h��S�ؐ6)c�m��*�	hC1��EU%m
mp�[��1k٘v2��s�w��f~t@���0Z���w��_��믑�;�S��t�G���d9,�1h�*�f���wP�b��3ٚ@��Dh��2�Ds�L@Ui�* ZkTn�lH��(<�g!	YR��Q)�D������>�':�睆p� H	���K�
�)�'�VZ7.��}�z�W�h�)'4M�c�[������Y�����=�j���_��K����o�;��������8<<���{���{Į��愫;�d�np��iʂ헿���s�q�����l�A!��Fp��Y�P�3��u�<zp��w�����ՖQ5fgg���c|tI��h��cO��;C�&�M���F
���q�<���r� �zt��I��E�Tt�݊��4��_�9G[7�}O�%�+V��zѢL��D""=��SV�S�L�s������,�kX�S�]�T�2x��h!�cjv]���bT1�)Fy��h���紽eZ%9��{�"���y�6�,u���kרON�̧�-)�^�������޻���?��po��hk����o���~�?�~��ho?��I9�A'�q��]r��,w|�P磟͒cD	^�'�<�H]���O�N�q/�;b]�g2���H	-|H�RBL��rx_������s�1�zL�J
r%�$ka����(�$۹���$I;�aR�� �G$蜅��˖���%��~A��MG	��8�h7�����{n � � r��4����T�!�N!��=H0wA�)#��qc��Q���O��O~�Df�¢�BGIk]��1w��fU#�q�ko�    IDATM߅Hヮ��}�e��%NG���u��]d4�e;�B�a��|�u��G�� 86i<��}�"׆��Y-W��1I��p���Sh��섾��4D�|�Q-^vT�g��U�999"��j9;a��3�cw2��)hۖ�k�F#�Ɉ��ш�d�~��-gH�#�e�Z��e4���-���G�����r���U0�
/C����w��k�ELƪ��<S���)�GR7Ghtf�Z��!�Jr]��2P�'�le�E�V߰qt�t�'<�����3�w�9����gT�l�ӂq�1*�x1g:��>��ǧh&�+7�����`׫���v`!�ď�X�ѡ�G②'��R+b#�8zAkd&�A�$x��v�������f���2I5[w���Zh������}XK�^2)x���⏆m0�e�r&�|���/�c���+����_y�?��;�|���������O���[o�Mx�m~�iKAq��[Wyn��Zp��?2�_'�v���n0)Ɇvڅ]���s�/�����Ʒ.��+�pα�-!v�����a9�QێL�BAg)2���ad0(��$����c:���+"
��9p�/���?������6u�	:��AKr)�c�J$19]��z�¶]-�H�$]ki�D	��aZ��q�T��EIVUD��������	ڐiq	{�T���%QK��F��5i4B���֚L'��-ҵt�%��O�����/}�Ljhz��Y��	��yݡt�t�C$*
��W\����������_b{c��N�<B�L&�H�5��5;�96#�5j<^Ŭ�+x��F��p�:hI��)����3]o����6=�F��4�s"8p6���b� <��L-|�N`=r)��XˀVIxFĀ�~P���󙢐�X$��2���m�s�F�R(��EϚ"*�F����1��
�w�cA�[ƹH��P���%����w������:Q$@��~2D�!t	$꩔	|�u�r"�Ƃ(�MESMx��_���������/Z����miږ"7
ں��x�h���wt�R`脣��՜���y�ۆ��;�µȘ�,��پu�2��nl�)$�Պ���xB�-��S&���=�09!2�Q��9����ΰ����X�՘�(�2bF�xzʝ�>��}���i�s�����x��<}s&�~fɲ�|t5�L0�0_.��f4��[��Q�a���Z|��='�N�ҫ"c����=�ôΰT�QI�ŋ���1�VH����(Rgpm��H�F	."uҧ��WJI�3	��阢�0E���Zl������8d%�����Wg�Ң��X�QW�ޑ��9*��U�bRe�E�Rg<���JJ��)��}!Y���"߽F��K>��g#��
���Lگ��9���f����h�T�*�m�<}�D(��Vq�.�[�G	�'�R��t��M�k�v�/
΃������ɫ\^���*U�M��W����������1��W��/�.ʍ���1���yp�����|�[_5[킝j§���A+��?�nV(�)��ń"B�:��/^��3^Δ���x�q(l���C��d��w��Dٱ���h2��`���W#J	]ۢ��]�(]:�)���jT��"��4*�����$Q�rJ���|����P��(5v����>µ5����`X�Vt��
����i��%�Yt1�9���Z�E��ְ�YL^�	ɼwآ`z�*�Wv�x���m0&Od�|H�{�n���{�AWsU\+X�? �"���[̛�B)��H/�nn��=�O�y�S����M��}��1�SD��^!�b�
��(�a�`kA�Q�.��?��sq����kG�Z�!$�����@@�@&�LB3	r� ���l�T �����c�����5NK��綧RD�(�ԆB����!5��a!�@�QB"e��P"${�(�2QV�^Lpْo(J��%���mL ��K|lM]^g	�:P_Eb��Q"}Έ�G�ŹA��8!�R���Vh1a�i�[/�����Q7� cO,��u���\\�t�E�HU�]��mR�$�m��)K�w���w���9[�ȴ�pt�>G�G�N��1���z�U^��_�4B2���@j�]�F׶�OJ��� ��^6x'P��xDI�,KDt�)1��'}�\ �sB��Q���Zy��6���o�_�u6�&�х��׃�%4����s��׶4�2X���MǢ�Q&c�W��	]O9"�l���=~��o�޸Mt�%�EA�y��_�"�O?�l6C���Q*}�L+:��s(����|�DWJQ]Y ��5�d2&���^���}�u�M2�E��=�gR�D��Ρd�P�q�<ǅ�����H�e�����u���W�����s/�v� �	ڌ�YN�-�1iNt�3��p|L������6��1���^RD��O纵�� �[��K{�$�o�?�{]y��=2���?~؂t V�	��~����x�v칐�� R�ܨ�����/����,�-~����w��x�?���~�O��?�Ώ~���n�b5��Wx�s���;?�'�Ɋ����Harz�by<���Y�ϺO�w�h��N�����&8�lL�޹�j9��}��f&9FY��"q��9����k;Z'�M&C�_ΰ�f4��S�[���W��ֳO�C'��gۖ�bF=[pvz���	���r���=��n~Jx���н�(�@���68Q¢�Co�Y�V{��l�
Wn�d��g����ƈ�yY���԰�(D��z�&ǟ|����}�O���8�4m��� �ݡ�?H<��ib��v��ՂO5yQ�ԫ������>�_uc������r[F)@&yg���װD���=>�._+k:ˇ�Kirf�ph��r��f�D��x6
:��	���:�%#���L5���H����]I��+I2^�8��.'������\�vRr�NL.�U#�L �F�#��+eƶ)@X���q�#� �$x}/�?2yzlL"#k����Q� )*�T�K�&K:��'�X��b������%�̓5�����Y����ҷ�鞽I��ABB�X(���C��cl�JR��rb��3���];T9v�r�Rv ��Hb�2H���H0�h4KOO/�}�w}�����ޞ�� 8]��������>�9��;��w�P�VΓ*H�KFR��55�� )δ���@L�Y���jPƀs�vEj<�H0!!S28�bw�`�2�,m0��o��l�X��lv�rc+R��y���iʍ!G�����%kgQB�B|
]��J����x@m<y���}'�W��������O��w|�sW�����9r�6�R�I�������>y����Z.���<�9BېHG�b[l(�kQ�R�%�ŋ�����A���e.ln3$�\�I=�i���Ȑq��@���u�$ӑ�+<2��JW��#�l�h��V����'�����ԝa���e���1�̐*�u�Olr�	��2��7�b�d8N��Ү*.�l�ki�{����?����e�E���_��K��+����ⲟ��n�+��O���������3w_�޽���W�޸E}��hk$�2�4�'��\=� �x��>%����:������<�	��	ޅx�?Yx�͋�������2�_g��ϳ�縻p��Kw�������H�?;>�}�S��_�����?{�ज़s�_���{�a��,^l1����E>�<r���࠳4��x��V��=������r�>v�o�&����#�<r'�� NYc�҃�R�hE���{�E�L�������7(�=J������@�O��'�6Z��6����]��~χ(68��q��ٻy�VB���C�SԚ�&M�tQ��9l�'[�<�0�褢��d�l�h�i��k;�siF�et�Y�>�s<]QqL��IЊ�Y1�ڡ�������V��jΓ�z�H��a0r���k/~�G�{�g���p��[��)Y�x=��.Dz�q�=���X����Y�˷�n֟�J}0���amnq��$�@�I,����K����P:!#�]��!���rq*k�@p��Ѕ O��#���<��P��s�t(!��;��E�)ВP$��b�U�RD_JC�xL"�2�tg��z=�8�]q�9��y �-D�'w�M�<
�߿^<.J��m(�9Y*I����Χ?C��Y�W��1��f]ͪi�F��`��6ض�5��S��=�l��9�1L���]�͒���xa(G9�@kjv�|�[n����ѐ�k�C����cO2n3�Ni����ٲ�jV�m�Q�#t�Dc�����-����p�Td��^a��%�Ҍ�#=S��bUa:Kj=�ݻ���*�f����.W��!ÍM�����f3��Υ; L�S�'SV��8��p��Q�iV�����v-��.b��I-��@���s��n���pgD�D�P^�7O��h%}�W �G��D1(Jƣ�(G�G��t�D�*��.˸�m���/}1�"M 1D�l)�)c:H�I�ԭݲ�H�"�$�b�I���۰������O����O�GA����?΅x�G(�����hB�{��P������[�K/Ӽ�2��-���mP��{ʚ�����#�^/'(��Vs�����g[�:��{�n�O6������U�"`I�� Q�����l^�'�3���K�o?��{���}�S�|����?�?��oy/r��^�p�]�fwz���1E�c�d�Z�)��Mq��9����7��C�V	�[�h�M|�ca!�J�����>[�66���SVՒ<�M_��SK��vΣ���iQB����%-�*jaI�ٮm��c��w�K����gZϙ蒨��P2�t��)�}��2�t����{��@H����,�S�U7a�^��4>Q�_`�s�$�|���>G{�L��a��,K��`1[�{�>��=���+���������2H��Rh���F�,�!�^��co�s��X��f�
��3��;���/�"n� +R��x�I�B8�T:f𮧐��B�d*��LX/�^�/寥,�?�-��%21!�	!�B��MuB�C�7:y�s�VR5���y��Z�T�J^�B�Q�I�L�\�XW��v�8E�#��T���N�'�
�Jk\��$R��A�Gۣe1d~0't)5J���3�
G�8�����������/�:�A���������.�Ӕ"���#Z��)43�i���)���%^��?c�l)�	z�E}#e��5.?�B'����Ӄ��ߙ�+a-����l��f�s��+6�C�|�����sWY�B@�2��˩Nzs��L�#�>�5�0I��ߥ13T�E���[/0��f���MV��h�����%��r������ӨA��j�B`����LIT*hWG��[��?�3d{���\��3� �jͥ�W�x�!�՜�_=�i:�N)�4�c�:Ҽ����;h��̧���rt�7���sWɛ�k�,�1�-,��Ӟ����i ��=���t�ι�/��ۣ�?�k�yI�j*��\�J>����K�}V�Os̨`����aNP�U��LR�!��S��G�@Z�4��C�jq²�Z����|��������ڿ���;B�տM��E��_�������]���7��M�0u��[iG����H�^�鸾����c>X���3�3����`��8��A@�7fY��ЋP�jCR�iHq�Nq$ٓ�9��s��g?Oy�a���'�iA~=�������?�>�K����|�9�&�~�2�����-�5�l3�[ж߂�S��}�d}qDT��_�DG9���<�ݡ��k����,sjΟ?�p��:���a�a��U]������^�U�1�.iɋ@���eF�f/�lڄ���Ҕ��&/��پ�v>�Y��yQ"�g�����̎���+/��hz�r��Z-�ꊍQ�v2Av�,������u�,6x:��?d�Ҕ��}\��W�򞧟%�2��N��pT�(ͭ7��>������댇��S^�J��a�HjA'[*9���Ŕ�W���'�'�����[�!��f�^�2�?���9&W��;�_��Ĺ|�M���0�|+�֒g��eT��J�%XBk��1�5��;�$>�ŏ�GF���+*Mlp"Z���6�Y�(2I�����ѡ鄦m:����Nuԟ���[��h�Qx2�Ht���2}HMc=�W8����Z0H�7��h}�_KE4Jr'-�%��8"��t@�[XMW�&����.0?<�:�"|A�5�8��ŷ�7 j	}���:뵶�zv�t*����s���w�@�*��HH|Ԥ������(��$L&�AB��B�]z�_��ԏ?��{��>�]�G��=g��]�x�U�jE=�s��]V��jŷ~�'����)(��9�~�7x��/���S�S�5�N�!
G5�b�!�%�f�%��!�Z�)3�b��-e�s��y�T�u�m8��ݿ���v���1�}�<�}�$Ys�F�p7�#�����Q��L&Q����	�������˘ʲ�������Pd9��c"�w�l�r�*�}�w����b��٧Я� ��[�@G�H=�p����O��c���+�>�s�{?�{�P�$�S:'��ޭ�T�#|۰�ګ�n�d��1[9�?�[�^��+�bgW��J�s����`F2�������:R��X�"2�L�54 Ü�wh��J��z��~ �������A����g�$����D�Ǜ��I�u����o?��9�+����)�=(��5�l��[����s��{&� &�:������%�ka������v�o����X�u�m�0��+�~o�=�K_y���������?�q]~��?�}���;�_{�������+7xx���,�~�[*�i;\��A�V3
n���`�v�[iVg��dh�o���ի���c�AʠAh���LʒE���mDV�����!E�PI����l]z����-�v%)1�p���ml��3��)˜@���[���/���-�w��o}��b�'P�5��c�m���XD��>�^&Dt�6�F��%��߿����o���_�ȳ�<���磓^��TBp��C�w��>����?�`���r��A#?y{��%�m�hrv�x���N�IN������k\�SV�)�_~���=C>~���~w��D���"|���N{����5���8A�.���{������� M��X�`"H�����e@`1A�X��4�Et~oUwUU1�lnI�(gPx��F�� �b���c¢��f��2J������)_�Ƞ�Ҥ=�y�<�ͤ�
�U�"�d1[���^#ORu�}gq�Ğ��eQ�@ʈ�_�N���[=�@���lcH��]�z�\�|<�� ��Б RMP!,*M�s0= �)�ѐ�.1�Lp��%M�l_��N$B �c��]n��*7o�A�6��կp���߿�l���;L���H�h�꜃�K�癧�VՊ�ʰ�����M]S�%i"���e�5��F9�ul^��p� �)j��]�R�y�,����ͻ(��L+�#�T�9A�[���uv����,f3��l_|��E��`����gwx��m���O��w?�+�	�R�f�bgs��v$JE�$��r��A�b[��}�!������Xۂ��	ʓ�9�Ʉa6�GGێ����SOp��C���$E����H�χ�Խ�{-��� ��8�R�Y_�3H(Z�ͺ#<�$����Q*����������6�<�B�Αz�ߛ%��F��E�Ք�5�i��*t�F<�������9�?0|LcHH�S���/y��3����$yBgR�	2�P���k\x�[��/~���?ã���7�4v��?����������7���c6ꑇQ��C{�r�#�Vk}���	���4�&�����шF&��N�8_0�|�nj2��BiA�DE2���t�z�%k���v�=��x�Y�q�]�ծx�d°j��~_H�N0�u�b>����LI6�c��GT���C0�    IDATx�#�d��ͪE�T�"�)�;���b��;.��_�*_{�E�u�).\����fr�Ѵޓ9ן|���1u�$�#E�T_w�Z��Eg�z�����l?�m�\#N�f��o����i�헸�SRn]����	�z��_���jE��$m���C�J
R_�������F�\��\@ɞ���e�J�q��j��v��xmdڟV�i�(�_7�u�s�����k:��R�giZ677�r~�Q�hǘ��)��r��"8MD/��e��b?#���~-�SE:�W�T|�A���O�u���$C���:�S�h>#t]u�����O�b5�Pz���'Z ��'��m��=@*5�����d�P�(���@��K���h�(I�ޠ�!�m�	����ژ� 1A��!i�-g$!��1��K\4���7ys:�`Y�4[��x����������J�봲���,����w�p���,��W�9�X,8>�RY�1u�iZ�
�ڒv��K��iIV��DB�f�4ï,ͪbvp�l��C�r�_�A�C�wv�f�|����dX9?>G�T��۬fKk0(���i�,s�<c��#}lٮ� :@ſ�D)�>��R����"稪���22�w��Dg4m�J3R��%L��G3��KI��h���.�`yᕛ���|����:l�����m�On�����F��FLKB���V�\����o`/^��P?��b�������{m/i��)*C��*��}&̛��ȣ	���-l��x�'�g�q��[;�HN��g{ԑҲ�O��H���[������ן��&�>^�g����_����7��|�������?���t~���l^�����f��mR�U+��tz�h <�3<;������S���G��}o�����dE�x�����&L%��#��h%N�k�r�F��֕�l�6�W���?F�ķ��+L��h3ДN2��t E�3�ɔ��L��*��UU�uJ�S��1�� 
��p��5��]	!�� �V+�$�,K���͛�mK�Z��1-B����<��O�[�3�*�WUE���J��6C&������=�m����[��)߳��kn�|Ǎ�dp�w_�L{�2��+���U�n�s�e�
i<}��O���11�KE����}�q�H���}�:3�ꆗ�k��5MF�Z;#鐬ږ��0> TJ���:�$��KLrA3�'������h�s&��ϿSj왾��}2��k��(�'ON�JB���?��8a*����(�숀Ht��ɘ�l�g�5�q���iE�?T����I�Ɇ���sgmnp��-���t,[C�(��h�k�XemGYB-,m�^�0������ʕ�d2�6�h,�[w�s��G��S/�Qs"�QQ�Y�X.vHF��-�H�t���֐����Ӵ�����8��,�wܹs��|�	R� ��"$!���f���'�%��$�뉓*�;�hW]ס��h����y��{�_ۛbL`<s�<+W{��ܸy��r�7�"�YE����s�����f�%:-p�Fc�u��u���t�(����g~嗩����~�<Oq.p6�ޭ���;�JR��	�x��K��Z#� K���s'�����NL:��Ht�@c�$8Kb*�t�S�|Ͽ�����D�M�gGv�����|v���U�XN�C'D|o:hZ֧�u���Y�9���;-S+��	Q��,p�q�$�H�P���K�\�K/���.���?���z<��|�����s�ů=9{�G��#.��4SJw*@sv< f8}�t�9�u8�O|����e��ҭ�8gY�j����E>�\iO)2$A��� tJ��hg��
���Γ�����^�G���dw�>h�\�x�Ӌ�"&Z`L�[뱶�mEElLg�#������ $��w�i��є��mn����#I�1 U`<����Tx��W�^ess{J8�i��j:��M4���O}���1�0}�k����]����v���s��9�/�Vc�Y�'r0&��Σ�@�5d.�1���u<�mL�d��$�D�vol�`���z4��)�O~c�X���?���i�w����Ⴚ�"�>ͰZ�!]@Iؘ���Ls�jư���!��p�li��9�������2�3}��=;�W��`T� >���%J�� ���U�H'�'%|�#�ޙHK2=)!I���ⵌ[�����v��;���>�'�A�t�b�1����lmOP8��+=�	�|�NI�Q[�(4��:�LRF�	�ł_�����O��C����ڳ�{��o����7h���e�̆QV8x���n�1A%h��F�g��I�e�	�9+,���'���s�&Q)��!�r���s�I�'���,G�%�zEY��7��SL�����$t6��J�U��P���&bP�px�2*3�D���X�c�xݳZ��{vwwi���`�u�����{l�7O����h���th��9��Q�߉X]��N�j������D3��/?�s�����:��t>c�l��fg��9�jH0T͌z~�sa�<�F�.��'y�Щ�dJ@�Syez��(G�2Z-�!M���]�x��|����A����7y\����oy����gvD{��2�m[$)g�4=o��V�y0ߏ��d#8���h�@h�C	h��h6.]Dd���>�]��<��߬k�O���S�������o�2<�0��p�c����d瘶���x���A5�}�-�����ι���������0L��� o0[�X6+�J#�FhI�T$i��RѸ��^Qd
�x>������-��\e����"���B4m��$�O}��4�~��!�,�K�B㥍���Gq{�5Zk��1�t�1��(c�k�b0�4�)"�lp�9�q�c䎠,�ႃ��+I6�`0�qG>�:jiQ)��1�o�&�/�ɽ=��N�ē\���ټ����_å��,�
�J�� ��i�$CwI�"U�� *� �$I�Fuo$c{-��ҠR
�o�ޝ�KI){��F%}��:p���tuK�to�ll�)U����2(2�e�d�P� Xy�Ga�����e����肃�(#��*X*)�"`� b�am��q�Jys9��3�D}z��~Ih�������}h;��4��I%#�x�D�{]�b���N�2
X�����.lnеG�{��&�QD�����Ķ%źRa=�x�h;_��~���#�t�7n����/���G7Ⱥ���$K�vxR��� K*�� 4�(�j�#�ə�e�I��:��$�����%�W��h8����%X��dJ����R�x��Xע�����h�Ӛ�8�"����tU�r6EiA>�����{L� MKQn�m��W3v����c��f�G#�4M�t:EG[7����Ɋ�s��욮n���	ΝԙD�1Q�Rͪk�VBp�U�k�|�ݽ1i��j
C��I���J� �i�"��mY��g����a\�����s����A%F���ld�x���4����%�>�]S����o��CB��{�������m�G(g�U��a�z�����z?��ݟ��'z����N{�'e� ��к�TD���&7P���O����ώ�>���_��O?�s����K��V��w1;s";�|Ҁw�g��?� �������M��e�"�5��M�Ʉn%��Å��
Z(z%����D����h�%�$���-�UC�=�L���Rg}Y��) TU��8gI2M���'P� ��c�����{+<B��xg1�=	�k T��H�ٌ��,��'��eU%5I��l�����Z���h:g�\⍣��f-��
������x�Cd8Q4U���=�7g��K�O���i���T�v���q�ݻ�����<�Ĥ�"(��ړr���DY�������2�)E-r���g���)�TQ�C��A`��� !��S�S�,Rx�2ckT0�R���t�y��r���� ӓ9)k����^N�ºL��u�[J�<-�N��k0\�i�JD.��!��� �´]Lx� IL(�R���(|d*�)�՗�טyR	!*�<���v�	�k���d�F;�xo9��WK�4��@X6����5˻{*a��e�����Cn�|c[RJ�3�yk-i��dB6�(��z5c�\�&��`m�.���'=` �	�f�*������� 8عx���dE��?�1�ʘ[k)$Z�D���dV�X��l��	��)�㺆��@�D��9Ǉ�8��yJ2(��4�����67���ES��j��i����f1_1��Z�����!��H���mɓ�,ф^�&IR�L	ї��r��ZDlnnrX-X�IT���	�x���4 7�t��b0*)�\ehW-��u-"Mq֜�O�5�\s +:D���kH��7�p�������G�����a�?z��/|�G�+��8�Gw�6�P �á΄�X�_�-�[��6�,�ln��4`���mm�,*׈L�)7v�r��Ǟ�&����x�'��SzP�<��X,��9�x<���q�=�['g�[����g?[RQJ��`�����?@H:��;:f�u\x�Q�=l?r��C�у!��sl]�D9��\�TU�����A��|��ۑi��&IB)tR�2�ԫ
�ml�Ȩ'���,�HӨ�B��^,���h�+�yG����'I�j��=����!m��US���EI���b@�=��n[�.r���FW�<g��ɾ�}Í7_�/�P\x�ݴ�6����3?ŧ��O����'�j-|��"ae:m<eg)�#35���,I:�m@�.3WQYd퐵��9Oj��$Ρ�E�-���V5�j�M���ب�^�4�]��jC�����jq���З�C�=T��S��<�xSa��d"�ܖˊ�u�6�-�$��[E�z~�>�8�`z�"s���{�I©��)F�4�y��E?�=D9}�iq�Cz�&�`N�F�̃|`���'&I�l����k��<XD������:#02G��yt��#���5�{�$#w�T(�޽��n�_����h)1�Ś/���"����#�&-G����P�)��E�;spPZ $��(2�DE��re���M���x�|>�_�/|己�c�\ $y���D�I��(�`e:/H���t��`Jh�i꺦m�jqdYF�e$e�C�eB�u;��3��BHA�J1Ǵ�a�XFIf�'�s�mn!�[Y����	6���>��l��\�A�XV/���8L�Ȋ��hv��-ZKD��	ɢ1,���*6�/HhZ��q=um��8ƞ5^;�Wѫ$�	Y������C��<��3������= 㱕��b4z��ܡ3�"I���g������y ��R��Ξd���nUB"�gK����&m6!\�#���?���z<���x�������w�FN!4�7��)� ߟ�Ύ������-`�u� ��~������F0���?z�]��wh�KFD��e˂�����x�5�$�!{Ë���oݥv���9V�(%pb�VK|p���$8S$�T"M����tBx�rx�DJ^�֔��h�d
���Ig�z�WD�q�Zᄥ�P�)�ΰ>���}�l� �,�9�b�C�nH;���NelT�]���M�[��w�ń��}���}��g�xt�����
�����9���vX2,6�v�2��\��p�j���Tm�v��+���i[J�XoJa�d�k��kw7V%�b�^K�.�%��`�2-s���y��,-<�(h���u$���Ƅ�R#�%�^btJ����j�2�;�J�y���AP���e���K�ӷނx-���EL(����A��Z��%�:�)I&�x�B� �BJ�V8���2�W ��}�>���]����ٚ�mp�~�kc�F�_���=�u�n�o-*YbE���S�[[���H~0�iвa<�hT���36�����l�QR�yU�1�m��
�5E���D�DY�n�߬d�2ԇ{\��M���H1�GHODŊ�����K�G��(��/}�U�r��h���`Y���	���z�R=G��.����r��Wؾr![d�$1��"`�9*#�̌�L
��bKx:��v���C�����+�.�"�k�jE]E5WI`4�(��9 ��PU�"��OVdg#�(�S4�����%� ���VL&���	i�S�:ʲe\gI��%t��l�sfob�;��m���4�@.4��F8r��uY'89c�W��@����ğ�����u��}���O���������W�G5��,�B���"�n]�Z�v5��H%$&�Tk胚�gu���@����cc��kEY�ll��\�o0.\{�����g��WAI԰�����[������7O{���O3ȷ��ק�D����kY�X�1%`چP������\.�f)%��1��}^����w=��o����$f���T��@��d���0ޱs���ߧkb֜x��f�m��e�$��0G R���|eo�`��t�	:�)���R�h���6����8i 8G��Fn�o1U��>�zv�%&d:�4-�i�����on�Ե����f��9׮l����O�c>P9������}̫��
m#��ݴ��4E�N6���`��,���y�V�;�D�����Q��u5��i�=Y[�:!{bCP�A��52L$f���RS�6�;�soQ�#���Y���!4�E�؇M��G�zf@ �C���7Xﱘ��E~^��ɾ��@��׷J!5�Iȃ=���f|=����{��5p�*�G�ǖ@X7�Ϯ���:�>=��_+�0�8:<doѡ�1uk�w��7K�L>Ax���k@'��[����}�Q����v�kȵ���HS1)���2�թ���"ୣi:�%�Y��8c4�Ŋ�����(��Hr���(vo�f�x�D��9�n:.^�̹�;��%"�����4-Y�P$�z���)N	^~�k��x�#c|ב)�c�ø��X�	��tm�o��m+ eY��:Q�1��L��4m��3-�{�aA�
%#�:)(u�v1Y��V$2|���̠4m�������P��E��Kq�f��Q2;O3��%XK�%�{�lm�II��x+��㮊��'{���h�[���RH:����K�H��襟z[p�#�p�Sa��wí��ٻI�K��7[����3C�@N����pV~d�,$i^0�l���������_{�UB+� G�-κ�yk�_�w:����F���0]I�B�}����j�LS|^D�����,KIE�pX�������<c�x�NI���ֈ��T�Omۖ���X,LFLjɷ��[մ�JK�AN�j�eRJT�o<�A:,#���Y�psª��V+�,�����ܤ�3D�W��X˂y�R/Ե�Ɇ���#��<-p�$���|���!�7^����!�O>��7q~�3�)������+��ٟ�¦b~�M���&�LF�Tp.d�[^���ي��q��K�'���|�vh��Z��ȅI�`2�y��Y��?�[Vci��AGH:FY�ְ`3aj�z]�qw�T�֊������0��@�*�"aT�d:�L�����:�^�%{%#O�h�v[U���$��tB��48�琱�.�Q�����@/�=E��t� ؘ\���6�X��F�h��$0�9j28�������@P9:OɆe�v�KB�Ո4Q�f�r����v�1�W�ie�E��B�A8�d8`Y�[G�����ZB᣼���i�����>�6

��[�uE���,:�C�>ŕ�cw��j.\��PD}�Q���߀i�Ya���A��8��8�s��xU"�hum��j�0�
�<�Z-q2tU�ЮI��1�P�%�Ʉ��!���:���3|���I�"�LiR%Y\���G�&�!	�! ���V��#ӄ�k1��x~@g��˒2O)�RI;;��*�ihWK�8�o���ƶu�F�w����`5z)���Yk�JS�l�q�����pr�!�g��?{���������W_��Я�    IDATT"���Z��wd��k�L_AY��#����u7q6��u�/ �?��[��$M�����b��|e�D��@��tݢ�@Dc�տ��,N��V��$Nˌ��n�ֿ��&(�ړޕ��n�x��tԘ' �b,�YT�3_.�[c�$�H�]}��l����\{�J�;GSU̧Ǵ�a��Ҙ�ί����1�������y�T������`qB0%�O{c�g�D}�kW���3O3���a�����.�g-NH��{h2�\�����&�f�]�$��g�z-K�;�ߛV���ՙ�M5Ð��,J#�l��#��X���l�������b|!��̈� ɒ)��(�l6[���RW:i���w�sN�&G�(j
U��޻��k��y���E�LmW�o~�ce�'X�V#�R�;c���ֻ\��M����$ڀ�
#4hI
�C�����5O�T��߂O�QBcTbR����\z�
;{{߹��:f�E�qi����'J��xĖ��,�>s�6�R�-�Wu�*%�\<ϥ�2�*Y���{�vf;���v�4IV*��q�(�IqrPM��C����(2�|ȍ7$r9�.E�0�R�{�Y���j!OIP�u��"8�ڠ&p��!3iq3��h�S�4�Q]�l�)jf�a��&W��!bK�ωG����Be'4,����#x��1j<b���)41f9\�PU~�0�;���S�%B$�q���.�
��d`�d_�xBl�"�B�DU��i�#S��5ͳ�z�t�ó/<K���WK�mI��H��a������򉫗y���i�?�m"fuG�u�mK)�A����PR�w=�(�^})� TU�;�hi�s�v͹�� ,�K����R��2'	"�@��J����"!���A��s��ք��r�eY2*!���VF0���(��]d°k��h٭jjS��C�0��yd�6E>dGJ)s���3׬޾��+����Rq�[8��6���t^�N������AJi�rҷk)eN�J�#3�CEkɩ��)�V�!�pԩ<���q�gH�S��=2����O@8N��+�8����qR(�.|:�S�H�;��a�S)e�{rCzQ8�p,W-��B��[���a��E>��O��H2P�&cB��K�߹�O�')�����?��6�������,N�ٳ��s'1�[������J)yꩧ��+�e:3�NI)��p.�j{۲Z�X��,�5.8����`qĢ]Q'�vl��x�8�d�/��>���������t숝da�������!8�W��$��6�P����C��(R�������0�c'�gIi �Lp���Z�T�����q��>�j�ؔ�"�e��(�%^��`$[Z`��s���
ڤ�w=�²��晗��ʳW1"G������v�T�����3�6��E�9c>A"����d�z#Z*J	c!��B�L�TRS)��b�o<�S����j�2��O)�b�p3<��o�����f��A�$�s��u�*M�A����]���SV!)z!�a�����Wx�%JU��3�e��e�x��{��s��e�����Y�<��i@��?_�4+VM��S��� 3/�R�� R����C��]�6��d4��Z��7HB���W�\aݬXV��e�-u=)D�ш�o��#̨b���M*�آ2�����y����w(�Y7}�x-���q��L���x���>EU����._���=����7n���=�mC׮�1P���hLQה�	øj��" y��)˂�e���m>��K\�x�g�{�w\��Cp�q1������f����
��۵$�Y����-�I�\���G�����Nn�h2�D�P���1?<b����\����G{���N��tB8t9jE��%��-p����s�:���E!����SE-gn�a��G<����!��Q���ܹ�
�=�M�-�C�����:����YW�G_�t!����+�Ć4�HF���'���]c]�v��z�	��������S���SO�QO���儽�/_a���;~��HU���,��ܹ}��k9��~}f6*�I*�x���̞���+P�!���{��킸�S�F�>X���m[�ݚ�r����4��dU֮�쩆��]t�E��������̯�*���7��Ã%����N��_�����?S����g�߸�(�kTI�Q���7�M�ș�C�%�R	'���Rt�l��l91��(�p�e��Gi&E�jE�R�DA�("h�e@%IIVA0�z�EV5I�L�b:�[r<?F�@%5[�&��}D����i{�ڙ\JI��X�F�SꈌL��.�@Ҋ����Dk}� J�|����t�	�H�I~ñ�h���=��zz�����_2RS�n�R���e��	�lK�5�S��Ԩ��XU�z�P5)�<�@Uɹ��ĝs�@m*��_b<��{��{)%�[V��o�����{w�RhC��O<Ͻ�#����`ow�T��G�IR!�B(�d$Pҹ�������QՌպŔ5��3������=�#xO���;,Yk��2Y�J�I�1��h���J��XL�B��((tE�S�\�z5ͅu<*���S��x!�(��U�'_�,/��27߻΍7�ٹG׬��2W�f��3� ����HRk}�1-W\�;ǳ/��'?�J���EӰxH�j)Q��*������}|pD�tB�w?��ʭX����y�&I�tK�!�Qx��8%�*!R���S�w����o��l����l��� rvH��<^��D�*�H5�HMs�k���:��fg�qS�m��-��0��_�������O#F�1�<��ܣ�����w�gf���G<8��!H!�_n^73�}J�F	x���}��;h��&�L+C�+v�\d���ڮ
EB�	Ѣ|kQ]K��~����;�v=�7G}������E>#pC��ͰcLCX�Ô��@L�J���^�;t�e������>Ef�N��٘I9���̵�*�x4�,v��E�6k��gy���H�����q���
��aM�)����������{�S��_���PG��[� /Je����C��s�?Dbv�8�lK��Dp�Ѷ!������~��6�ʀ��^B@�DE6��B����h,M�!*Vѳ�4�1�st!)�	.�v��%��I��tm�-S�6/��P�+-)��*I���J��$Jm�ƪ�r�R&H�6�ƅ��^����>����5��l��T����B���;b�x�<ۣ+,���7��8�	��H�%Vk05Z	�]�@._�����SO�޿úk�x�"?��W�����Em���\ƶ��#���o�����G����w�x��ݛ�� �IF�d@ˁ�հ>�x�qYv��bIGĭ�W�a��y�qN{�!�syk1\�h�]Ǩ�h��#CYU��˳n�18B���a6��������Q�1�~�KvϝG̶�����X�O|���6�0�!:ۨ�^@���^���_�o����~���1��Fk���!F�d�ߜ�m�lMx�Os��S��98'E��+O��5����< �:Ѵ����(Ƴ	tkV�CM�y�/���߸Υ�P)4�|�fpi�qQ�$�"��U��ݦ�:|���;��.��'
Bd��	We�N=����=���^<Q�KD���o�x
���9���mXϏu���[���(�1��G���6�K=��G!��G�;[�6_o��f���u��6�5"C���IK��)6�!%�(�I���S)%�Z\��H��z�߼�Xo��aqD1��w���Z���Պ�耛ￏp���ۼ�X�>8�?���<F&�xaμ�S?Ƽ���e�xg�&F������moq��E�j�12��bgo�3�)5;�	!$�r6��Q�"oڮ�=�i�J��&����~己��K��4�Ǟ�{�nr�O���/��ӻ��m����	2jt�Y������8F�-.Y�����y�3&5�'n�-QE�(z�7=�:�5�ҢG��P���(��خS���g��֓�b�KvzM�J6���#h\"z��з	5*
�T�A&�N���W���]��e�(BD��A������kA��K�i�6Q�O!�Q:᝜��L��:m �3�I�,�c��@z�3�N옫�&
��tz�s綰�!HK�z�N�lb�,y`<��ra�y�>`�ko����K?�)w���`TWL�5�{�����Y�.�0��}�%�z�-�޻K�#��C�n�%�f�t�5):��֑��c��L��l�bB�w����g<�e��HJb�ʆ=U���i����lG�,B)�sL�S��{�.{]�Ӹ�'	�Rdӭ~}H�,��E%���������{|������8�dV/���޲8ڧ9>fq�w?�Flzl=�R]�)R�j�ل(%m�捓�� ��K���(�U��(����L�S���|�����r�CtE&�^I���S�ݽ��~���y���]c����kJ$�*�aE��,#�;W�>��?�|��:���(��(�{1�@��8��e��ZR�B��4��G� �@�$�����P�5���`��O����_�H�cy�/�k�,�"�jRג�.B)OBh2��I����'�μT"�� �'���ov$��S�{�R��hL���!}-<���%.�[��ɘ��<u�&�x����]����4�9��1v���L�$n}���:yj�A�	�
A��͜���z�o;�	�[#u���I�Mi�H��n����yܢ�[�;��#v�1w��w�GKo@��G�W���}�Z���N��׊}+دz�H����z�X�{4c�m�(]P3Fs��0�F�8C%s�Bni��S�Vd��)rZ� �,Y��L�ٜ�͜~���9�<%��TD��8�B�EV4�#JJ�q��_׸(h{h{��!E�?�X�ƱS��[���j�״�Y)��d�KK���R.�jcw":@���X'�� �Ȣ��X��B�f�e;:��Q8����u�	b:�0�r~H)��@�8h�!)��&���!�1�lF�2.�%�Y��,��Q�e6w	�4wԅ�����h��.����������i��Ã�s/��x���+f�mb��Gk1��E:�t|�us�����/�5݇2�-j��ܰKJUH�,�4����25e	���d���O�8���hW���1ٮ�}g������[�����*��RaXU�I5��U�Ry"ms�Ȃʲ")���[�����z�M��ѹ���)~��Ȗ�?�i^��Kh�A�e���� �"S��r����������׈ﾅ<��tVrW�M 
�����q驫e���#T]�h-��Fnm�G�f/����%v��2�
�v�%m��z���K)E��n�jG�Y����5eQ�n%&Oo3��*�H�^��RN7��;��U�b�F����!��k��X�����������GhDC[�luAɨ�{&����)K�G�)U&�
��bD:��#D��4x[?2?�B�L�w�"�ii�~Ľ7��勯���#�\;�7�����0�$�ǽN�W�L��Y������O�+���G�]fq=�Z��F�.F&!b�	�ːOZ�(����V���(��Dt�<2E���C���Ȩ����Έ�l�3zcJ.��ۆ��H�)]��&{��Q.���&�6|Je���Ώ�jXG� Mv�rC��R��Q���[�v�V������#1�q�ж��H�`�ŗ8�S_�;���H9�Ex�J�UAun?�HL۱=!��&	|9�5�T�����\�g��Id�p����L�M�(�0F����Ѓ�MR�$�6$z��}��AnȔ�S���7�ˎ6���(5^ff����J�Ͽ���(9Q"��mFz*E���Z�TVڴ}�h�q{a�����#ųS�n�0EF�-�^�ф��h`�
��gU�v#D>R|<b�����f�(�M����!�%E��0$�%hC�Кp-���dٙ%F�#v��QB�z7�,g)�����ki�9}��N�h��4�5�slᐽ����!��9���P�\�JϹsS��E{����1�R�X̉2�J޿�~f�Fx�h�kL�p�1�F/<γv=N�TB%�G�6�^���Մ��uM��NPVn�ޖ�S?�9.>��}C�%��L�Lt}�[�9�����9���-�v�u��|ݢRI%%�?�].�s�Z)��1��0N�P�h�1�j�����S��>��.]b2�h���M�������oQBP�&��R$D�F���)I��F�D͉�u�^"��xI)Q)�c �����,��鎗��+���v���*ʓ�(�jyƱ6"E�`��;a�A3��]h����D���B�@����ٹ���{י^|��D�O��"�sl�(]#�v7�a������F�Ǟ���Ʌ���f��3�dc�#m��CR�:P���J��TW��s��將Zw�(�i��u���7k�vM�)@���=޶���J���&:�^wL:˴�(#9J��*���z�:��
���E��6Kn���ж�q'r��낲�b��/Z!i�����EᛎJ�H���r�3���/���+���L˚>��z.|�%���}��(g"@H]dmvL�I�L���n`V�l�ъ���S�غ�ו9���њq�)��i)ddRVh�IS�2BJ�ݚ�%:�C""QB����+�$d�R�$�FU�BPhC
�-rRH�@�y#��5��1�M"EO�Z�
�LV��DRh��!C�d���!��k*ΐ�b�GG�j�%v�����J���_����!�����@>�Db��D�  ���L���q]���T�7-���q�E��T�g�F�t6 �DK3H�����|�b9'������tK�*Ҕ׶H�0���0m$"
��$�{�*y�����В��^��/~��zε�|�\�hZ�T��'���KL9a4Ҝ�p����.9~m�A�A�Ct4�9�:�0� �FW���K�[���u������s�+�8��5;�Iv�#�m�@��+l�7���M�姮B��:�F)�l<Fc�5#Q0���c\*�&[�7���wL6aY�VXk	Gy5?<by<'��&S�x��+Fӂ�H�=�DDԈ�s��čOʣ�s�#:d;�AĞI!i<��Ï^����o�)���=�� �l��c��^�Ǽ�Ɍ^q�l��Q�?�D2�(��0�"Ks��׸Yl����Po]���;��ꗏ�8��r<���2����!�<�1|?�����l>��OlX�b��|��2���j1x��l_����B�-�s1J�dYX$֒�[\��|O��������;bJDr�\�o��o��}�qY���â���Kl��">b�-O��D�e4Z	�utM���!B�TƠu�v����QL�3B(�KT�=F[�N���|�B���6o���PNvx�g����/�*C���,"E��r��׾����<x�5��PF���6�CuI��O��8_s�y��t�3+�d����qag�3�u>/}�O�YX�!aà��XM�������[&���t���4t���a���@���h����b���l�Z�䬃B��\��i��S��z\�Dm ���$��b�yͼ��E����E�,U+�x���r��#��|H��9�0ϥ#>A�Erm�m�������d��a-4o��;\�ݺ������v�r21ѯ[�G��5m��뗜߾�Jo����5D\L¦��$Re���#�LY!�f��.Q͒Ż�eK���>|�5�b�*h�&cjS#ܼN���΅�H�����！xp�2���FCr,D�4���u�-�[��i����׮��̳l?��h�#fWs��v��]�Ժh-&	���?u�������]D9\�7%֭��I����C�GFjD��uL�d�HR��}�b��[�2��"
O�lom����[���/o|��װ�c��Ϡ�!�D�̇@)���)QQd���=Jk����w��<�{��xH��w�#�    IDAT��c���!��� �g�C��*ns���	t� T�>�y1!bN��"�F���!�aqL{��ϼ̭�_{���r�GR�n���o�������j�먢��t���~8RJ��'C�O��/�?)�<7���g�C��)w\""��yt��a���R�T��$>)\���"�G1�����l�����{�����]l����^��$&C�[���O��Or�ӟ�u���Q@�
?huuRx����UubX��B�Pj��i��Nq)Q��JY�k��1*C��ڰ]*>z�u��`����x��a}n��AE�����w�����f�'_g�<ŸB���Qf�ܤ��O��|n�ə�#���w�AF\�x���E���H))J�w�;>;�� ���ږ�לT�G�'� -41%�%�(P-�.Q�g��8��ad����z����^S�]���� 7e5B�>�u--�F��h��6ЯIm$���	���cA�$�=�Hg�1!�D��KST�2����	E�Q�ݣ��C_��b��%�Nb"�DYWhJ
� �xG�9��R"BOX���>���'"�Ii�2�T��<���%��w�F�r��TZ��)��L��V��F�5kT��]˞�)�,����� (@׿+^�������a2�H	Z!�>��,üS��"�T�v]�D��&x @=�[d���]ү��$��B�e}p��7^㎂ŻX�V4�%��=B��AnH�Z��c�Z��&�޿���me�Ibm�ͣ����QDZrr�B0O��떬o^�^�1���m��Ǯ�l�mEQ�&��s��XOg޹���w�Ƿ)�=	Y.u���9�a3����9�D2�i�g�*9����e�x���o~�Ŝ�t	���x�
��E�(j���So�!�t6�� [q�+������(K<à?:�;�9��O=)�����~�ս�/}�����qt��/����^��ަ�s�1H�,	y�~7���I��0�_��G.8��M�Jn�R��}����=����$����"&�2٢�� d��R;?�l�C�&��f�yQ��1@�"�D�}�͘����^`��A��Ĭ�hb��j�6� ��0.+|���0��!JJ�$#�FgǬ�B�i}���P輩)#223����L�@�e�#��mn��Wx��AH�ňX�ip��0��J�P#M#�%�J���G��7B��w��t������4Rh���$._bww��G7�mK�?l&z/Xv=���DJ�!�eB`m��ђ���]�H��Y��L�����CH��g/�(��1w���Ɖ���/>�D��� �\��a�P��5��l�Z�0X6��>Qr��I�	<�:˨��������"&F���7��h��qʨΚ}��>	";����"����Ѕar�2/������
���m!�V�f3�>��k;�v0\2]d;j-]�a�CEA!MC���)QI�⊱.�M�?O%8���7 v�2)��&*��pNYh
i�%�ɨ[:ee��v�BjCR#D���-J<��=��ضa�{J�'8K�p��{�;����T����b�\�>��]��E@:G�-B&b��-��E���e��W�M�(����9R�H
-�)���#��X�"���5�C�@)"���I�W�,ǽ�n$�Ai&�FW0��j�Hx�("��e�>���Z��o)52ETTt&Q���{��������g�����M)�<����R�:�	ZA�x�Ǔ&�t���cr��h�!761�F��a!I!��cL$��4��(����[_�*/���q�����w�~�/_}�s+�����_����U�}n��iW���Ȋ�z=����Z���I���!+�����c�<���$IJ!�$GL�Ƭ�����`���1��L��Nn)!�Bh�wB���CG��1e�����dA%RDnܡT�^怔��Ϸ����ڟ~�TMKY�(FctU1�ؚL�@�n��{���TEI�s��2Y�(]����8�q�Ĕ*�,K�.y����u��I:_W���Ï�3 �HL1\0�%�"�z�����A$�P��"^��N��yL�|t1ȹNeb'P����A����M�sKb1ƙ	�����Vs�n��=MX�=��Zg������o8O�DP^@�n�����|���ۄ.}KH��vV}���L�I�{\%��(Ifi�����R�6`���#Lh��˶A��Ai0�M,۞�)3QX�����8
R�X������^��>^`���N�I菓�B&Ɲ^���ײ��		��NU�l?�	���g���@�YvvvH)�3��x���t�9v��Y�	6s�����&�	�6�����	1��6���>1�%+	�Q=u$�X��s�l0T.W��
�G�Xg�b)�����3FQ#��b�]�$����W���'�6��)#jta�,�����`w��:�b�d�#��.��ۄ���)�X��������z�;^!G#�hD5M��dK%��2�Bj���B�H��A���icr���	�G�|��HH$)�.Q��Y��:9N����N�c�#,�p����Ql��K�ʮ�J��:`��^�����_�׏����������W��{@$�11z���Ա3�{�>��^zx����c$Iy�m��24�S�B���ֺ`=_�ܼ�������~���ʿ}u=�x����_{�/���ۯ~���%�sp�.#`�9����_I�}��o����*}�������B���O��ic>���HG�#{J�"n�'���:���S$�P�P�@O FE��6��(�&��B�Q���!��J���b��(*������{t�c�LiC`>d;��)QAe4��4�$v0"idQ`L�G�)G�U�ָ�	t� 56zj����l2�ЮH

�M���rV��hJ��!+��J������P��:����N�6��3�II�q�Y�WJ�<�03-��m�)��{t�r�����sj�����N�.)tQ�Er��O�2�	�GHM�����M�޹]��RcYܠO�#]�XuEv���jVQ�@):���Ao��#^��Ȣu�U�������Z���D� �M�E�b�\#(�˒�2Z$�Yۆ����.B��^|����/R�%���s�7(�{"R�q�̣����H����Փs�4��k;�VG�;>�l�c��%�SX�a��GO��D��Ӗ��D'pn4��-](1�����&�1ED���y���?��[�d�+*�����3��Wiz�YZV��)(M�ozJY�|��vk	2B��$zg�uE�K�	;)�Mp���l/�һH:��
a*:�U@(�)k�P�w.����n��6Z@߷��s�YM]���vuL�h��_g��T�eϑ]$̦{�$q��4�,�~��7� C�!��0��s��\��UV$�@a;G�AW��P :	zo�B�9`J�Y
��4�c�{u�q=��9��ЮW�.��H�6��Ld�3r�C�i��v��V���7^��)�.~�Q�)%����{oQ=��	A'�aԗ!��#�3(��?t�+��"'���3��
 hQ$�#�v����!X��%��_���k{����߯����y�s?�C)�_��_��������/}�4�����{�d��ւ�;�*r�W���$b� ��!@`󁦔B)E8q��	u�aC�ܩ�$�I}b��;�S"J1��-BH�n4�$[ll򉖂� %�gP1�#�^�&������[` �HTT�Xd�U�
������5�����b�#R'�XJD�I"�ݚ�Ĵ�̒�!
tU�UI�Ȉx�s)�(�5Cg\	|ʤ�@���j��Dq��(\�0l֬(�O �@���O\T%�o誀��Bj���cL������D���b ���sQ�I t$DO|&� &%tH@���I��(�) X�a�Ɔ8� 
E��_�DlZ�y�;���Y"��I>GҦ�)���4r�3/?��g.�n�$�]�T�B�\�y��w�HD-����>���mM]U�՘n��s�gb�.jR��?���L8�0�B�l_ܡ��al;^���ؕ����78��C�[#d5������ɼ��]�Y����"ZiR��AJ���z�}��-�����G��+�p]��v��]՘j��Pe�4E�l����0,�1{��R#L�-�J+M�I��VqM��αՂ3#l4,Zϋr��)dt;��O_����9�D��(LI�Y�HuY��H��0eAY��tx[�𪪧6�#��\1V��Vjɹ�ĩ��s��)}�a�t�p|�lg���6���j��Q�fg4cO��c�%�H�튭^P�%�E�`~D���������2�Zz�h����~�Wy�^!h���Q����]ߒfT�h��:$oE�V��R!�@��(J����ح����17R�_r!��j��9O�Hj��hH&P,3jp0�l���������O�����h��I��?x~���`�M��yX��JlL���Y��y	$�ޓl���RD&|���I�Y�	� �ʄ��}B��Ќs,�>����6����/~�������o���7���~���Ɗ��w���o�O���������2��o�o��.���(	)K�|�]�V��=e+n
��u�o��:�?;�}��;=��0)�3��S���G�]�5�ٸ�[<S@R�䇟.�q�amP�Mo)�9�?�����Y.�d���"B!�<2w�z���~y�s�G#�QH�����)e����g��?��&jx�C_?Г�%�=��:yl|���>W���Y���Ӣ͏��ʹ"o<9�XCȡ:y�(3�r�E�}��(H>P��o��x�����m:נ:O%$�Z��/�1ۓv��]9� �
���O�$$�L��B���!�G���k��&]���o��{�~�[\c�$�ш�9yu����2>�|o���CE1�xB(��g#\oQ)�"^��;��U�!�re��b��
50⅒�����^�9:s\0��a�[D���xL��(��y�^3���x�u��_�3���w�mM�ܞ2.R�x�Q�ʊJ+��հ�.)��dݕ��5j����=EY⃅�4^#�k����v��w��{���{f�Ҥ��7�6r2�ٔu�2�H՘5��������y�-�y������,wy۬�g��8�%S�Bm�6˖���$��?AA� �#:!0p;N"ñX��I�c���/#g���{���r�鮪/TUwu�s��p������]]��W߾8���b�0���G�52_�ܹ�uC�Z_�Jw}�ю�̈�x{���8��ay���g��a�� ��ީγ87�.���ln�ke6�3[,q!�k��@gQ+X������zCC�����,<�B��2�{,��ZRZ͵��o=��_�}�G�<���?\GGz�2���֯Э�#���.���%OSt�$^��Y�zez��<z#�k������L��p	1���_N��k����_d�:������/��G��?����S��{���������_����_��=�?󧾛���I�/�F�̦��xCln`LM�M�\c����[���=��4L�=�qz��(�0��g.�����`$Ĝ�!��o!8��˥Q�͂Y@Gk�a����B�<��!66KXT�\c`��㖫��n������ֵ�̙U��s�ڙW������LR۲�����\4Cd�+��ξ�iPe�5N������;v�U���(Nc+>%a"�"ɽ�8j��XW\u0v��7hO��u�;.Q�w's���7��5�f��%��������Nc�=U�˟��o�b����T��p~����֛���+��U��6��}dJ�6�ާ�/���I�x������jźuxױhj��5;�õGHw��5Ǵ1�}�tG��� $����x��+� �*������K�G����yM5ߣn���k7���α~��Yp�->�0嚝�r�C�-��ei�m8���W����@D���l1��愝���+*�qZ��G��O�ʗ���ڀ�Hŗu�g�u�-�4��%�#�]�5�H�!`�C}���5�7�f3;3\�@��=<&\~���En���pr���7���O���N�l��N0��m�qG]74�K�����y�ut�5^�f9�T1�2�n�0AY�9��p�_��DF���J��P�YH��l����o<��_R՟������f��������gYqmձ[-8:>�Y�!���,��T@*��i6)�"�>G,�j�� �4����c���/qk��=x��/����Wx�G~���У<�ů}����폞���^z�߬��W���_����~�S���'>�_��?�];���_��^��u�-mbԥ:�)B�253�F���-��d#n;�1���9�|�0f'Ɩ���4�	��@�"ģ  }�b!��#���>W�S�D?���P�a(���8kSÛ,����T('��������!�7<w��y��3˺[Q�E칮���Ab��	.a�?�`^�p���(T��6�TN_�S���wʦ�³i��D�[ i�hj5��D�Mo�'W��>Fޠ�$�L���6l8��&�28��z�17[��.X��N�5�������GQ����gb��R�2v��q�yc�z�	���!�W��HU�i�Q�)�S�|�g�N��� �]��C������g��G��U�0�@� !��'H�Ӵ�e�Ν�x�����}�=� �9a8x�2�~��\:ڰ0�\S�l;�ٚ�7ܨf�\��~f]�����M�p�v��rC3(R�EMfhk��X����J��ڰ�Σ�.��#�|���:u�c�D���2c�X�«�^Z�:�ɚ�d΍uMwp3�onn���}f\�j���\k��J���^����x�e�IK+�1��RU�ƂG:�7��`حgԪ���f�ˈc�㼏�9�68�gO�~�tw��8*�V5�W{�(�l�\���:�=�����~��g��1�b���������[6�F	f��;r�6%s+Q8֬�����Ķ�ek�*ֱϵscN����ƒ"�������oK�6;�ivgx�|���_�շ����?Ȫ}��߸��o��'>�w�],.]����1��_��������;��/|�^�~��;���ٟ�I��n��-����.����q�#vL(�hC��0!�i��B�1ҧw��G�Ɯ&D�+��-�ަI�Wi���)&���&�J�'�\>٢%�A�$��U�j�ͺ������sƻ5�nt4����qW�]���Q�$�XJ��ޱ�@Y� �'O ��bҜ'��j���~�S@����Qj���!��B^b�!�XK���˟Q�ռ4���P�|<��PG5���i�t�[��h�x��U�_��]��]�*hvf8\PDb]��c���="�\�9fK_��'D�'k�=�O��
����\��;�%ө���6�=hXASp�sQ�&�Tc7�Lw�o���,�&(N,�mp"8�ؕ��*�X.���푃�~aB�̮��@u�#c���Џ��3?��[�vkv��x�
a����.��lf�vp��3n��r��{�a����?�ct�<����_�lZΝ��4ur�t�.Vt�k��%}l|�Ժ��i�A�85�͌�߰r���ªC���j6]|V�d4
)�$��ڠ�fwQs�>��l1#����9�Y����w��������O3{��	t��gT��O������X��T������A���c\��-UP��!���7���j�T�\�Y6걳�"��9�L"��e�Jp��x�sZ�"�Oڬ�"�g!5�y�!�2�������_�ko������?����m���G�v���?�kO�����o��]�Wp����W�;s6W��=|~8���-Ir���u����5�l�I�P��������޼��1,��C7-��U�����\��G��{y�v^���[����폾��U��1�z�o������o���>���r߽��?��̌r�my�[č�<C�    IDAT+7�n0?�����zx���ַ�Ӑ�z# jc�P�Al��,M܅�z ��̌�Z�6��߯��gg��?S�|���=��@uV��N�"<i�2�o���uX����hd��<�G/�a�(���teV[.�-yX�M���{aŲ���X��m����M��=9��݄>b��:|d>�0�m{�͕2��{�V�KM�9k�9�'��$�1R�8��N�|!�����
kj\P|�XUf�$��J����GG��[�1�5�U���W�����H4��QC�s��x�,[r��$AC�G'3D��B]UQ�433\ ��Aƴ&k�Ӯ��=����ht��sYjye��]�1S��]�oŌ#�$�R�"M�$J�r�B!�-A�5�T{\;�G~�G����p�u��	��~n\����'���C��=�)�Z����a�oن����d������Ƚw�ҋ��@N�h;�nS!p>�[O�!
C&Rv	qO*oq.��R�8�QpA	��Z�hlWl��a�;�+u�"z��y��_A{���3�O��������w|��y�{>����/j���*o��$W�����k/������ɟ�><��g_fvpL[՜��?�]|���"'{sNB�l'W���\�nW����>�%�o�9W7x�Ҟ�^3�u��G��ؚJ<���L�R�B�Bߒ�S�L�]2���9�To>ϋ��������z�_���K�w����k�����>����s_b��rmp�Ҟ�+%T���Yil�W��,t'�(5�*�?��J�[���%�~��$�&�+\F��,�b�x�<oo�Y�\�7�S���^9��+or�3������A��v�K�}w�ރ��_]`��13��~���_�ڕ+<��3�j�~�P-fX�,ｋ�Zn�z�X�[0jSQ[��1'�g���yd����˷�to�q��\����,�R���I��U;��˙HHBYa��ɦ}�S�DIm(�4�lC4�q��QLҌ"̼*ZW�Mǥ�S��1�̪�������8�e4J�Q�L=���2�[�`���cs�Դ�͂R��T�ضO0�<���Ef��汉ztO�*�H�0;�*С��`U�R��)����q�48	8���2׀�]t��@!��
h�胲����Z_0�A�c�֝���$
�#r.�*�mn���6�l꧟~wʢR�x��c#��I\� 2؜.�7Ifz��6���=T04�,I����.�|��Ǹ���'�䩓[p~�>�<�����G��S�@^ycg��;�﻾�����B5cs눯�Ư���~� ��Œ�۰�,��t0�b��$+�@l&�����y�N#�M����<>cFl,;+5<�2E|tZ6�Qvvfl��,t��M`v��<�3?���pp�%���"��%��� ����������_a������x������
Ǖ�����ٜ���K�3�fE=�,4
Tn�Os����?�/��GϿ�Nepj�lx�݂v��"TZ��
��1KL̈́~���{)�
'�����֋O�n7uy|���?�ο��^8�����o>|㛟�'���o���.��X�^��#E����es�����e�Ō���AS��39Ɗ�ʂ~��>kV%�U4�����l�Ys��?�ԭ뜰Dd�|�CX�G�s���B�	Xw����Y��u*S3�wYԻ�}Wò�����+��	��M��Y��`��XíЁ1��NzSGE�q���ؘ7�⃦�;���4�$�����1�i�ۙ��̿�Y�ҋ��~���*�4l�1=�+d�(��������^� ��S�f�*5�	O��ر�l��M�ٔ��Y�[{��EM"i�Vb��rZ۶�^��H�T.�_
O����v;��6&T�/��O3$b4}n�������U��ʫ�57c�u����-�V4f��@c*@�����;ܷ�������M�J'�]b��Zb��b�þ<t����2�<����ƺ�-c+����X��)]�@W<����h�^l����])!���J����F<J��Ēh:hmX�Q36VpP<&vy��&0�y����������+Fx�o��(7^{��ц���7n�p�{���L�8�O��/}�ç����,w�d���[S�P��j �Xk��-~EB�sŅ�l���u�Pi���&^j�r��G�
���`mEmRbkb��5T��t�������#�p�e���/�����Ks��>�?�=�����'��!��!��\z�a�}�}�u�eړ[�U3t�q����.?���`�G�:dy��؏s�w}��8D6Q*�AfP��U��:
���:Î�@�,����+E�e�Ն�A�������n����������~�+��K��=|��绎O!����o�ܸ�G���_��;����k�2�8ٟ��ќ��a��u�YE���(`e>�������0�>���m������9ʾ"��L���8IS�� Uo�F�ZΥ�t��+��Ҷ-��8�jkh��\�u���8��u�J�xU��.� ����]��1�X,�K�7#bD��f*!�UT[���x�����Yi��?;�di_M�th�Pj$1��x��opY��h��x��O�RRSh���-�A%k�a���i8gKs��������F�gJ���&���l��6�����sQN�F}��],����3n
G���1�F�ɹ�:T�lf��f�0�������G�n25��Z`�y��L!ܕ������۴�SV�,��2�TN$��6g��W�&�6��(U�N�� RWt��E�P����]2�N���a�9:���?�����M���]'ت�s�u�:iڱڈI�Wt�>���E%�)r�2b`��;,�/V��[����n�X�<�S���8;��������n��YI�,�EcI�bO{Qct����1�s`�&xG��ص��'0���q�8\��wQ_?b��K|�ſO]yv�5��s��#�w}�ø�*_��K���o���1��K48ZjnՖs)�^��>�S�ulk	���5f�QS���Y݀�
�Dw�HLÊM�t�~�T�f���"(5G͌��$4��+��g>�	�]n~�Y�|�+���c�q`��囼�~�ko��c?��8?_p����݊�n��гYV쮏y囿�l��V�=��?��{.V�����gv���tu��tq�jwL��0�
5���Ұ]�E$�c%|�qT������\��ھX��9��n�d���/�g��[�?������?�������?�=?��)�p����ˏ�����W����_�+�\��z��ۗ9\�X�̙�C]�R[wb�1�����eo Bt�ZS�s�-5s�[DԦsiS����gN4+��g�{6QN?ￏ��$�O�ڼ�ſs5��t��~�
v�xR�ۅĔ�M���<dҢ4ϩd��d�/�;k�g�����dj��ZaW�GT_СZ�y�^I�c������Шa�����»�x~���;X�b�:!����p��kgi;G���x�!�y��}�K'�F�ŕ|�h���9���]��4��ɹc��=�g�ܗ_���,��W����^�\�j�[6�Q��ž��ǭ�uYA���Fs7ոÜ�.?7����S!)=t곑K&��=z'�K?/w;�?k�2��F���_���!��e�;d����wq�\pН�g1�kg��&��T��>�?����c\�r�Ǿ�x�	������g?��?�4���u�RuZ�k�o�t�\Bp�]�cS[W4�ڝ�J�Ҫm8��nS�Y�`7�cj�/wؿuH}n�����U��u�m����j���>b�س<��G9��\?>�2v��t/�=����n�]��i���]�O}�g?�;t��\�/	��;�[/le	.��y��o��< [����c�6'kB稟��E=>��������?�;_\S}2T�?���v޼~�G �rk�ߺ�;9~�l�~������O~�.t7�㯾oS�;*_�A�Q,���V�(����Zlw���M��v�+k�@ʗ=�~"g ��=Z�u�U���r��}��&��,�5i����8Z���g�?�ۺDS
�	��m�L��ސ�@�B�X���D�TAc�D�~�}U.��G���(��3� &��^b@� �h����kϾ��z{����7������t��W1�)��1��c�S<�����Z}���?��c��L�|�yq;�L�1�����Rt�
I�Ph!��gaI�j���w��/:ش��O-������Gm+5m�q��tNA�^�3�v�!��&R��_w
/����6�J����ǲ���gb� ���Ӗg���:iSP^������,h�U3N�]��Ϲx�.��9�n�ij�[aW�RR��A���?���{8Ys�{��]�Np�w!�1�+��\���r'�	�Sk�>��235�V=jbS)<m���fͷ���І51��;;@�:�v�y׻�͍�6�t�f���"��j<��[��Y.]���|��+�egv�N�ci-]�Q���;����y�s��:��_�%���������l��i8٬b�U�mZ\�Q�Cu�o��7��4,B�A�jEc�Z����/r���q�=��λ?���Z��Ȧ��#�9Uex�2�/��Md}L�Z6+Vo^#�N�'�>�b�J��0uCf��Y[YY�@����=�t��UeM<��N����&�������kl�v3���]	�12
��*��0�q�V��T���ʜ��1��q���N4���O`;1���s��ޏ���5��z�}�*���ޟ�^Mj��؉H�z��MǋϽ��6�l�g�
���%�}��VR�)�k���<FIoOȷZ+�7Cszg<x���=q��������h����a�qZ���qk�9�\��_@l�[Ѷ����<�肀Ԑ|����9�����:R����~�;�=�,V��-�M�o�pu�;<�*R�^���`;kجZZq4��f���i6-3�\_\�qd+�Պ��}v/,y��ț_��wp����C����>>�S�Ͽ}��z�]���ê�=��:��A������֛��O�i���竩,����c��9�{�ON��;a��s!,�x�[1�k�[#'G���!T�*��.M8���.�Vp�Y�������!v܆�>�;��O���XB`u|B2��B-��/�,E[�w4��2ݤ��|<
6Ů����A���6�>K3�1?��bo�P���c�9�p����O�hW��x,�����K4�i�x�������%"ɥ��7!��n�������1��~+�?҃Оx����~�mf��f�61�@�/R�_6�T&�G{�.����	C��.nwm�b�]K٦-������Sߏ��~����M~����#���7��<�B+ۄ���a;I�l��ZW���;�x�M�I9�;�]'����T&�"�����L� �l�ʰI�jz���ꅳ~���'�܆cF8�m����߉]
���:Ì� �5��x�Ȉ�{T<�������2�,�(���N	�جM������$��*Ov	�Q��6�2^�>���ΐ�Bs�B��Ti��������3�,<�(���������fya�p���/p�R������a�ܓ_b�ݝo����s<�����`�y��?�ݏ>�+�>����9�`��3��,��,7�k��sB�8<>a��1���շ_�m�`�R�l5��
�9�*��{�=� �T���T��	���:��+�[�\I����!�7N+e��J=W����G������	��	�����_���u��n�NN�>Ԇ��i�#lZ�U��Z�h�k
Sz/�����n��G+Z�>�TR�L�uR��^����o'+և��)�%f[�Ϫ�Jb��
hE���߀�Bc+¦P0�&?v�����4c���C�g����F���D�)�G�Z�ۀ�䠝�Q��MʹASy��S�1���}B ��MV�r#s����uM5q�)!�#���Ҝ��,p�9�&�|����k!��_�� 
�'l�C�^ɀ�cg��[0y����K����J��6uC5��c�������3���s�X����C��ޤ��jf�������]Fb��Ts?�ɗ{Q�m���řȵ��A����ɵ%Y8�XN_�����9���c�|��6�ؓuX���|��MQ45\�$2X䌎m}ڮ�G|W�Ǚ�m��iky�߮PQϩ5b�LI��g<�c<oy=Q��h�G53\������g��[�p�����������������o���]<��?��������xϣ�g>���^��+�nR�[��.�W���0��去�į[���:�E���{A�v��`�7�Y��A[vfU3Cv�S��/�x��.0��.��ជ��3���q��Wq���.��朻x����!;�oۖ;���|���,�ޒ>�����g8�l�%�c�5B%U�|0�(�BSմ�bV}�.Ֆk�`~[�����&YՔxN\JH�`��t���kX�����VAL��hq�l�X�'hL�^b!7,�9�s�Ԑ,*�%2�^�˚|��K&��F�d<��{!��+ж����24����cm�}�r��i�,�����r`�9s�߮�wXSj2��( ����%�ٖ2�MЉ?��}��&u��d3k��Z|����u������O�@!�'E��1�3J�4XkY�6m������_J+���7�B��~��r�6�ߓ���tn��8K;��{�瓹:	�r@��X�9�)~a:�@�f�<�	���g����۬��]�TU��y蔡1O,b�{]�d���W����L7[ 㪶���5��6{� ��P��o�z'\�v�?�|��~��[�1�C����\��S��������h��:��#GW��7�������C��]<�������>b�9s�p|�/��'���/aև�ΝG�!�dPaٵ�F�+�X��9��
�v8}z� ���%�+K]��u͆�����56o���?µ�9���#"\z�A����޸A+;�������︈�k����2������>��G���'�����ϸ��	�obv�f��X�!��QI�$MZl��X݆q�z�y�{&8���]mV,R)���EUqA݆��kQ�upxϩE�"����ǢNjll�k*p���a$e� � ��l��ޘ�W�`�����"&Z��}U�)ˈ�{]��6:�S�q�å�}A�����jRJTD�U�oF >��ՀļޘGI�@��~�(�R�)�k�~gA�4beM?���b�Z����ٌ"���W.^�7�ȂX�ܨ�{9�-Z���=m͠X}�.�&Zk����Gd��e��s�@u	������o)����H�)�ֿ?�MO3�&��z߉1�W��'�6����ͤb�P�%��`sj�/��fM~xf��x&c�����&|�	�
����#h�p�]G%��]Ƃ���h�1��1�~2v"�Us�q���!J�&W~_^F��l��p����q�7��?3�W��5�Ն�>�\k�|��~��>���Si�;|�g?���Žz��kG���Ǚ�s�=rΟcg�����|�����o�:{W^��ތ���9�g*""�v]���u�����U6�U�v`6�)"����^[����3��}�<����G~��~?����9>���}
��*�����A��nÅG䑟�A��y��ޢڽ�ރqt�U���_�����s����s י�e�������fV��|��[�rۚ��6�W�߾��hϛ0��7����
*�5M��pX��Um����q8צj��n����xUASC׍�ۧ�Nב�BHe��
 a���"��V\�:���U6��F�F~�/h4M��g
^#cp�Mҗ���5��c$��ƭ\%��Q����}u����sx�����4�&�AH��Z���F��ܘ�(~�\�  � �(~}�&��j�
Ԅ�Xa0y��'��|��,��y𪊥";�R�����KG�ؚPZ+��ҷ���YM=�� e湪im�    IDAT�T��7i�B��נx�}��lƚU�)A(��K*��������lR]c��m]�ԲP��U������0&���0��D�OOL��[C�f2����*���V�&uRցFc;f��M�R���C*�M ����*�:��Ezq�Qi��Z�=�o�1Ǘ����w���}ã!X3Y �=7B��eq�����Q�S~-�/�HAi����@���V����w%�Na�0�=-��8�X�A������gY�s/M��Q���_��o�z�*���c^���98x��`ynɝ�]�~����WX����}N\`o��3G�] ��)E!!��Z�v��.����&�gvR�T��O条�w�ݚ��cg3�|�˼��+T�~��G���`�K/��淾��?����#��S	�s�v�6��^i�չ4�x��M��Cf�+=�����-���KTf��*�ex�ͬ��Qb�
����<M��}�scA���h���r���4$�Z��X� �����M]<A1�4�T�9��E�Q%6����Y�;���H�&+K��R�j$���<jt3m*�=��n�bqi���Ȑ�zBU�=�W�0b���i�L2aOJ�V��"}�:52|��S�`��@#1H�Q4�2 @�b�����RN�d���1c�5�䃍"`zF#�5� g�!tUH؈���H*���|D�w��(=��t��M���^���cF�^ (��ɻ��2�PX�B��ҝ?5���9�{�oqH����"���
!b����%��[��x{�e`@�=�(?=$s� Q@��`J���R�H�gt(�-Ƃj�ed����&�	�P�� ���gl�šBYY�4���h�.�̏��qʊX��N�=�����w�l俳��@gT���Ѩ�����M�<����¯U�y�f��̰��٭�NY=��|���c���w���D������'4	��\�]Z�N��1�J��l	�.��h
H�î����ڷ��k���q,ko��@�����<d���'<�/�)�wpb�u���"���kC�����x��	3S�O�ys�	kzM��x=&1��E�:�H����CbZi�m��v���1+F�|��3��%�ޟ��!)�f�#y�[!��넀	C��L�!/m����Vz�\��'++�7e֓�4lа�ާ����	GVV����O���_!5��%_)Z�N�ʔ n3y[,� ��O�El�4D�O6������P�M�G��������^���Ӱ.�[��H֞3���g$w=N�&}���E���;���$�ng��U����	�9�4�0��52��"_Gf�3ĶK
�l;�����NA�Ɣ�X�q/)5�K灢�6Z��e�.�����N0=mXlQ!~j�^�.e@#&�Y���;Ef���t���t����3��N�T���p�4�d����1;j#�F�	��1S��do�ύ�!"T�eU�᾽s����"�5޵���V��-��c����Κ�'7�2�OI5>΂�"S�~rՕ��#Vg4��=k�9��}�7^���%�k1T�c�f5��p���W>�.�F����kkt�8~����nc1jX�V�1t�b�ABSLW��`vw�1/�02N/��Y��=�3Rƛ�+B�s�yD���3㌡ms�r�r�ɥZ(_
Cφt�F�FWrt�+�O�p s���`���c��QD8�ç�I���6Byzqф���#�f�9��D�Y3���ء�����w҈�kĄ2�J�L�R��L�0��T:�����-=��ACLI��n�LK�0F��V��,�N>g�Xv�������ݡd<2��I=��N�ߪɌ�z,��/�L-p�L`>��R�LU����sg5���</�w����=i5Q�ġaM���K�GN��d��%�9�i?�,�x��2� �CWŬ)�r�~k�p���6�U�ƘΫ�|DS'4fP\�k]zZ��E[+.x�󄠈�(ڶ� �T@�!�dRo7Ufs����:�Z:�p�1����h��:h�NJW��=)jx?dMd<<K �p{�3��0u�ߴ���yݰ�X�;6��1�?8��9�+��p.���jF���*�@�zj�p1t�ۖY���.�Y��U[>�=yOR
\ĵ0:?�ّ����S��r�����O�)1���a�2����~^K�9(a���w�d!f2F
Ƌy$idYk�/Mz��3�(�yQ������h<?�6�ƹZ�D�1���0e��"`��I����ArĢ�Bl�� {��|�Wa�T���%�`B�dp��>���D�C��ˠ�DA"�2�3�5�g&sJ�D����KEv��o��֚��C��vbn�G\
�Qd+����O�f �s�b^CTm�2��DoG��{��.q�����pl�HOi�e��s���ِ��G�ǿGU[&�����z�H�s=`"�p�O��R��X�ςS	��{�d�x�>�8ߛfA�Zd˾�{r���e?���F��� �� �!8%t�؋cP�����Fb���)��m�x��1���1��[cM�x0.v����k+�R�b��`��w[5�w�n��Rճx�9Z�Ҿ8*Yҭ��i�[���b��{�<�x�l\`#�z��S)TM��u�i{�$@F�%��ٌ�_�V@�R�Aŏ�Fz#��\�R�֭��o)?��%�.�H�˔���XQ�0��K�[U�7�9Ee�A�FO?DݗZ\p�5��Q�/Si��Jm<��l���8^X�U�y��$儐�Rz�*Z�)��K�K��n��!z�Ǉ��jBxP��V�`��I3<ҿ��$-��]��S
 z�RP^b�3�^H:�A����e��Ж��"ogE0�4=b庡\m޳����$�H*x�`Y�4ǲ�_�_?�X����0��IjM9�GH���h�3��Or���/a<��m�?��gae����Y�Ϧ��t�OQ�}�^:Cy�4�G�Lw����#����șk�odd�,��b�H�-�����{7� !��K��2->�h�~~�Cq� �|�}��y��IP%u4hXQ����X�k]s|�f��1X��Q+X���4g�j�BKO�{ׇ�-��m�~�����v� f�<�8+�X|J��.�Jf��'��c
m�=ud�jT��5f�Xa�Y@[�8Ϭipm�.(k�6��Ta�SPX�"k�y��Hnn=��dV�g]Kr����m0�O����mV�OΈa���l�FW����
NB��K��MD���X��0%��[A�%�a��v80��\���6�e۵����	�mFH��g$PU��/+���@|ۗ�b�B1Q�C��~��k.e �iN95CDFf�Ba��� ����N�����|
F��;�7�,M�3��p����0E��~�BH���
"B�b�V�ߗ�8����� 2Lb8�cS2�%���4n�O��ʈ9L���8|fF�gig�]j��[�If�!�(h!Ȍ�ʼf��;���Rw+a�s.�sa���/a�)�;Y����`q��� {s��&H�-�$�#�Y����q��Y����0�*�~|�Da�F�:#�S$���X��(�;���14H��]��ǊPױZZG��.	e�bd.�����H1*?�<�,�����"W^uUc���t]
�6�Z��������n�Sefp����t��*j*o�@�:lUG˦�x�w�JnQҴg��/[i�>�5��y5���T�J>oy>_f���L=��\��4�fz�9���|��%�(���>�0TJ�o9�ؼY��sZ T�@�}֥Ij�p�A��>̩�Mk��Y{F��U�4����:�sTs�|�z����m?Ŧ~�is�S��� �E4�����i�HL(1��\��U�!@L� z}*Ѐ�9��,b����gF�#/��'��'��Be�s2��ZO�UO��0sGm��3қ��n�~�������� ����t΢%����4������宋}[��&��s[��Ո�B`H��a>��x���Ê��D��f^SD`Y�=nL4u�6&��NϹ_�����WP��K�C���VN7%�J!�l���m����~���������A`6����fk]�)^R[�ڮ%��������6T	��-xPk�eZ�^'>Vz���8������г��xou�a4�
� �V��77Y�`B�ewg�r|t���kq�JY���Z ްZ�]UQ��f���kDR�ƺ����]ÆM���:��Vf�Y���Fi!d(ʔ�z%�Z)]��aVfٜ��Fgۯ�
B!��P�ҋ^P��l4Dc/,����ɋ�.�� Fcd��04�|�pT"��/�����Ny�@�n�63�����h��� �{�m0���a6��*k�Y�����hN�y�u�!�9UUE��E$�d�U�O$�<_IE�M��4rd�q�!־D;:�!H*���-5�L��*Y=��̀:DY柝��p��\��ѻ�H�
!�گ���EQ�Ǜ�H 56z�;�(@��bоpR�2�9���7�$��Pi��M�п`N!d�H"#�AL���-����_]b%V+�mb � P�A��,tq1Gׄ����[��/<���/�W���Ѿ�V���}�t���)d�F���B%Ub\!�c��EWָ��FgN��2�ȁ����UrF���'!���Yr{谦��3���hza8h�t�^���ArC+�F��$!:�h)�yo�Ƹo$%�i�^��
�&e�	���Z�,�7�4M�+R�h��sD�������D�Q�����V=�q11��w�fFc���	�E�}��EN
�Z޳��g͢��h �
�`����,�;lB��#.�r��
3q��/��v�u�5ӵ��u���>�:�=��¦�S!le(�X�o{��ު�
L��J�Fx$���~/�w���)z��9m~����̛z�ؒ6��0�%58Ӵ�$,w�%��.�d~T��I4k���M'_JP�Mg=sZkʗ$�,���RD����G�N&�����]Ef��i�4��nǐ�3D4g�%o[ԦB�|"!j��w���/?��,�T��*h%���!ˡ���� E0X�W�^G��G'�aq�SM�$���A(`��P��5�^�<w=��M�͇4�,��;龕5�<^pmJ3`���j+��{!�qPG���fl��:�/gp�.����{�����݈���,h�7��S��3l%�i�K�������CcƱ�C^M��M�%�Tf&$7:������Y�>�����(@��n�1�!�>'٨�AP!`��@�'�#Dn����Bgd0��ۑ&:��1!�7��ˠ�T,

)'����cA5.l�Y��BJ=�#�`�C��-R���\���!���ͮ�����A]H�؀�"���2ۊ.gސ�F�3�ĺ	�z�Q��rAzd(F�n�pk'�y�d�DV*���:��8CF�U�m�'��FlLq��P�3M��fd�^y��1�1i�9�j����2�0"1�Lu6���o����n��U�����E�C61���3b%�> �$F��T>k-M�P'��b�/���)b�sf葐��l6.���_�
ǟ:���9/��E�����62q/��1C�aS̫��|S��Ϗք����ZY?�YϜzm�B8�Vy4��ؿC1RE��hT�%ٰ̏�#�%��3/�y�gf�X&U&�{�s�=4U��[��'����g��J,e��Ks�a�~�ʐr��a�UD�杪�eKSI�EHn�`C��V�`���O�������Ĉ�r���q6���T�K�;6Yx�Thj�@B�j�0�5f�ы�"=����T����O��;UM�ȸo��<=1����oo��"�!�c��s�?�O�s�f��ZX�b5�E�_������Ć�N�@�1�`L5��4Df�^0�k
���(�7���#@K�+8�t�h�a:4��/�ջ1�L��S��3TcS��,M�@9u�ƌ|�1K�:"��¸(�=NB{!0�3(� ^A�'øw]����,��׿���g�"X6�W�X���J@����x[%��N"�����w�̉�R���AN����i�
Ӌ���Pr6�DI�Gٳ���`�!�L-����Ĺ@�����5��ȁE��B�hp�&Ǐ�c7�`�+�T ��wnI7��J�"���ǃ͠� �*�i��͒s�ҳ(pCKI���g=(���N��5��T��Ϝ�P���>��L���"@F��%d�B��b��>�T����q�����	�DCtW`��0Ehs�>1��R�H�u$�7U�����1D�M���e����X�\&��KsL��ʢ�\-*�,��
�(��S���|F`�O���A�s���lnV������ُ�����f����0P�qK�����G�!ƚ��b��Г����ݦg��2��>�C5
�Cy��
�`e(Ϡ�8�k'[�����I:��3�}_�9��~��t,�|*�L�	tܕ2�n��[���)22��6�qJ�ma��&��TXp�PC$�����C�~��OT�:ҟ,@ga���q��l�0I?Mɦ؂�w������H��Xb�4������ݣ���
� �E�~�^� `� - �b�g����23��^3#�@�̮G�H>S���~�yxxH��9�>r��Z9�l����F� <�{?�q =F
=���Ǜ�WkIn�	I�ɉNptJɴ�G~�J:N��A��ч��D\�g[M	C��Ci��' Ɍ�>��)ұF�L�mx��~�(�����G,�F�����PV����m|��;�/�Tn�ÈtOR�ٟ'��/�ww�w��f�g�ObD9�ݣ�����"Q6�\�&��cg�>�-�����\t�[��|TA�a@��Ȋ{��+!����(Z_�W�4(�E:5�O��2�a`ꒃ{�a;�3:�+�h�Jk��!(�d�u�^��P �NC���F�C�P��TN�[�u�4�<lR���A؁��v:8�b�����?:T�����:uB���/��҇�x��e)g+�Ɯ1%?�	���q�12+���[�e�p�}� ��n<s��ιI	�f<h�' ���].���}�lY��N�Hɐ�S�n�������݆^�_<�?�s��� b�KN|v��(�]�4KY�Cp?�	�8)ƾ'/ǃ���qp����~�#���ID ��o��^V^'���2�:�vD|t@�?��?������w�}Jɔ��6Fz�����{�g�����(������@����F�|�Y;胛Ï9��qY�X(1A�M?��Kc��؜1V4KE➤��!�nl����Fqsn?�۩(?QPE����u���8�z��[W ?��Ǎ�-���	6�����Ά��C? ��6��P#�<�cd�4�YP��@��J82#��CWS9yCы�H�Rt�">����B���"	��!�$vO����$��vT�r6ҽ��{`�v�^)�����Z��ܧ����PPN�@뼆���u��AQ��b�
,�c�:@�����rms�'rM�D�v�9~~-��#:]̨G���Vܙ�~}��f����o�*P�av@���r4�#����2�7+Rv���x�l�����6�1?�	�`|�pK� [��y �AY��.��^���B��l��g	Tr>k�JW
��@�L��5&Ip����Gg�8����)'{>��N�$�>����60��71��A�ފ ���ݭ7�z?�_��Cp���.(� �<xS$�`��DuD�D4�)Mo�|M'䉱�C�����Ä	���`M���N��A�?�>�}�R>�@�"�piG���=�Mon�Λa��u�'}1}4��oc^�� �Au:1�����c\�ł^��;j+�L	�Sk>�2�����'���]�^��\�v�\`l���I��ʾd�7p�`qc��Z�C�?������?�����A�ܙ�)�P�s�"BN1v���9�q���g��{w�)*�y���`��%�����"#    IDAT�b�7�cYc����\���Z��:TfosmF�G��;��	�)�hZ���X$�{'Fg]S���XO�΋�X��m�BUL�Z���C�6�ۣ��;4�_��Mr�;C���Z)���z���}D6\�	�[u�� ��O9p�UZ���e��X[c��t��Ck�U����gaMS��p��} E�j�V1瓃�������!0�Lc9Y�aahü��D`c|���t��pL�{3�������{�?Z�
gc.���=^9gl��ǩ���٩d����dm���i���6�	���·��F�p(�RR3��%Zv��B���3^�c�V���g��	i�sla+�f�4�����B�Cyx��gG"r����+p��
��g-5Q��d:W��h���P=4���*W�Ίa����A[��I�#��|�E�4���d!'n��)l�(ሰ�H��}�
px�.�A�"L�$����Պ�*l��R"Y��o� S��6á�@5�\����gҫ�=z�6�/����U���X �T���2dV�2�z�42�Kmw��(��ƿے&"rV�s
H\�a���-׏���va8��_t2�T��hvD�e�1��6u�Fn{Ygs�O�y�;|NE���A	�p}Oj�2��8�j$R_0'k�j������{#��We�>:.KM�;�f�Z�n��,���k]>�he!�>:1�q?E�L�|l��"����}��s�~6�M&��:���_mNʇ����s����QN�=V��f��]����g��FQ�+���t�ugԶ�Ef�	�BG�ָ ���l9���,_3/V��u33(g�.$�Nu�:uBa�����z�"As�^py~������X^כ�o)�(!U���UpSE��;���?���_q��P�H����ޚ5q���=�C� g{�.���p�Ƈh�n��r�6�v��@����w���i�"w+c��*���ؼ��`�*	_�]�MF�y���B��4���(z��)1�r��0 wj��ٯ&�.��3��Q���hI�`�i3�jl>!c�����յ�����4 K���_�J�G�j�~;�	�l(�U��q8�����Y�8ٳz�U�>�ʡ����p��p� H��*���tj�KA��@i$O�$F<��lƲ����Xf)�(���M0���h��)��!�g0"����4�ӈ6�)3��ض���Zt7X�ε��X�L��/��0�)_ 0&�vw�|�[kPG���`�Rpt���r(hK�֡��PkG�^@ʨ�Y�^�Q����W2�2;U,[���j�ɮ]�E���N^ƌ��T�ԫ�������!�I�nN��j��Q~��{��ooo�r�t��$ ��+)e���lA���`x��O���c����Z̰}�b��e LYwCU��I)y���>˶���l$��ɷqm��ө�t�L�3;�����"~�vAfF�t`�# 1���Am ���*�w"�*A3c+�#)�$8�qX̩'����:G�3���lz��H
\K�1�J��>D�l$6}%`�^q ��Ղ�C � ��ݣ�V�`�d��G��ߐP�
y��A<����c{2h9�hḲ&�v!�����;�\�u�S6������n��V�� g�@ZOx�����Ě�$?zj�<��!e/wA�~�Q��.1>N�����\Ԁ2�v��q�D>ϗ&t- �+F??(�8�8p͑�%�].˦ѱ ����(r�h�9JN#�!-�B�+xx��LeJnP�3TGe�òIeB�s浢<� p�M9�C"�B�H'A��  �w��Tf�'�P�w�ȕ�@a�մq��g.ڌZM�(��yc7���9X���g�5��`.h�Z���y�cs�\�NPZ����m��"��ldґ]PI�/!>�����`{t�8�����6	�ŮM���FG۱�l��"�I@�� b<��V=�4�pGC�&F���$�Y�!0�TȤ����
�^���&���$��"@r	Z%�9,�w�趔�.v�
8É�@�
�����D�h�&0�[;�.��k�è[�CL��jx�X�o6y�6�V�^�!V� #sf2��{�`��@*	�a��99=/��ש臭�ަ�Q8�#Y"�Q =Z}���*�z�5g^�uE⧓=P%�6�D�T�G:ɜ��5� p6���	��v2��ُ�%!���dG�zJ����044��[F/%�����@��߃�D���f�lrNh!>A�˚�0t��{�����|=~xr9'��W3�M�F('�1O{k�D8�������VG�ތs�A�zN�֙à\=����/_Qoo�r�P�М3���e��#3:�gv뺘��̐G.~�Hs��ilV��"�ɠ�1����b/	{���duƦB����N�PG���o�Y޸Fk1��T�/ش�{������� �;�G ?z�xߡ9!-KŖ�Y0U97���6�׵��$2)T@,�(��J�"e�#I�Y��lh�LU���d�>��V�
�^��{�j������{��ٝ��@�&"��n�}Y��O ��:��b���8Zw¥d����q���M	G���[�5�NC�� �n�V��[��b��^�� m��^�|}��<-#w�X���GN���9�X�5��G��ԇ���f�b�`�p�H:
1n��%h��l䒑��`�ޱm ���������㨠��!ӅA�lG����Rg�&�u܉G�s�&Pe�DeΚBXQR#�*�RL_�h�u?EFw�՜�!���wCcΨc������B6P�����>]+���߷;>�'�7@ƳF
��>WiiC[fJf���y3�Y�q%�c�u�y���6?;v�ws�������m۠��j7��BT�j�2�<�(�[-@6�ު9�p�.�� ����6Ќ3�{�S�_��Bnr���+�
T�w��GC����A�O/S Y�Ŝ�sB.N@�2�-v8���)����+^��YT����u�!�W�{G�&��H���j�ʶL���/l^JD`�ٴ��d)��5͉�m�^6#��9Oeu���Σ��z�U�* Sg��|�޽��u�Bn#"�H1�� ˵�I\�Z�wp����Q�;�10��Ύ��3�_=��~<w��p�9��� ��n���Q���C�⠜6��D@�D0b�w'&�1��w8�S
�r���m������R,��c<��N��Z+SJ`'���=�Y�L��o�����'\�i��v�U��S��̜��t�&���rI(ŌZ��R����;�6�l���;R!���I���P�/��V �޲�$#�u�@O�		�u\K���97碃����tttb2C�͉�"h ��!?mH^����� �]J~o�����2(w(
%�PTgAuhjv�DC�k) ��(?�5L�]�v�5�ۻ�:"����L@ڐ2� � �#�֠�S��HJDF�+�{�^v�wyC��?_���w�ү��5$O� ���*c���ɾ)%��X���� �@ɢ{��gL_�U��q@�5��~&�1��&�m]W��h�91��:���D82���J�8c��9c��i���Yp�c}ϒ�����5��Qn����8�������l.���� ��{Ux�+�5���y���K��<,\�z�����z_9g(�P�Skr����Z;�����p����uG���V�s��_�b9����ʞ/��}x�� I�?��0�Q��/8����L��d9Ե�	�Q�+Z�=���mТ��a6Q�L�P�K�ɍ\�y��is �����ȼf#���\U������k�L�e���0DF��vsqc.�`{�(���B1�T��J��aV��2J�b�VX-q"Oi�N��E���(G9"2�Bch��a��K�`z��[+���w"�*.x�$s*�o߀���!طY>5	Bs.A>L5'�vk���5QR�y�d9��8�D�mk�9�JwuI�咱��g�qTGE�Q;n���H_Q6[W��g���7ʟ��;�"ؙ�f�'d9�a7��L��}���v�X��U�%���B�q���w�
�:��զ�(�v'�zΓ��������}����;n������ �6��/��ۗ/x~~�P�///��n(\Pr6TQ+������1��r[�W;��0�5���?��qX9|ƥ0����E�`K/�d���-�i4{�eS�/�Xh6���Q�*Q�T5��UG$�[3\1�P�H����Y����Υ2�0�<��z3'	0Ni"HsG��^Z����0H��������bj�W��W��H�v�#���h{yƏ����ϸ��,t��vC�x���o����m�a�U��'N����-|}ư��b�(-?7�n�����ٍ�Y˗��4kMil�x�ox��7%��>dF�jz�2h��A2��O�n���6G�t�l�s�h�����R2Ja䒐[���1��@)������E�hn�uR⠎EDoa3����F�$�b�*<��G��ƺ�W1������	����f]������8�0c:a1�����g7�v���Q�DD����q��ĐK���E��˩X͵�~����h7���[�cYg16aD�݁.��:h����@�'�u�B��-�7�lų9���n�:�R%���^1�p��/GɎ�@�WD�_�������M��M��j�wH�͊Z#�d��ao�%���ĸ�\������d0�/�����]QE�(8:�W�@m�A��`f( �[~;����[��w2%#��\��g1�Ug�'��Rv�ځ����h6Ykuf��W�gTvZ����nJ��� ��F��:�O�Ƿ��@����������o)���ߍ@!�����$i�t�HA���MMc:��>Ά17���ׁ(�噶3j���x��}τ�cYe��`:S�v�k�����i�
fsJb�[`1���w̃v�˲n���J� � �Y���?����X�·���3ǻ����@����6���Z)%Nx�W����Ox��dN���ϟ^��� R��j�qqB���BŏX�"!�������,,j��S��o����߳�r���㘌���夰���K�{+���^EJ<{|Ƥ���F��c<BW�~�������w�����O��N��<�7c���;�NH��h1*�TŚ�IN��U�ci3
�ذ�ߠ�"
F�-w��̖�����&�D��fx�F0c�5F�f�n J9	.��@�f����^"4���L(P���C%-hM^����[�a��d�����5(wO�P��% �4Fr�  g����i��ס8�|"2�5����a/���H�`Pݚ�(��P6�N���SA~@1AdN�H�.�l� r�������"$��J����5rZ��w�nw�	 &\�N�ׄk�z���p=!����u�!kC)����j�{�3ZKP}��zE*-�^}CD�`�ɿ�V�;23JI�vX������P��t ��+f�S�Q����r��׆�8F��֚�&��e��9�6$�u~�E�W��8䔰�+jo�v{�O��������3������xzyƧOW��rb|���H/��A�w''t@��8�8#s��w?ܷ���X��G����ZW���*\/� ���(�� �^��)��6�hDg'$ C���6��0�jG���>�K���qHH��#ؘy�H���������P��v�.U�6��w�m"9��l�"�1*8���!�������ҹ 2�S�������xz����;�\
��`ˤcߪZ�E�3&�(�����c ա���'�_e�I��V���8NY���&�/�����8�o�}@���������o�921�x���	e��j�ߵ�*p��E��K����׋�6���p=e4# J�w�1���'t��l�]/&�::l�r=��܉z�v�=�4�E�q�^�o�VI ? ��v&�LF����lHM��|a�#J}8�<���~U%h�Z��U#A�LD������A��P��Mi���*�k6]u�Б��ӎ^j��1�cԲ�Ch	�c��q�g=w��ɟc# ή�.�y6d��<Kyqv�Q{��W'����wU�5��mL=m�lH�-׆���������W��V���|��d{��8�dK���;�`?,��@�-F���x��'\.WH���Ў�[���7����>�e�������Yyuh6r���r��pI�Vz�q���|��u0[�u�M�Hd���hM��ml����L�D����;c]p;���m�� �t�z���v�ض�?����~����>%�O�=��@;^���=v����Pu���=�R���R�;�����r��6�7���[���>�3$
��E��- �l���X��zX�s�p�Ww�u��9��+T�M(���8E��L��_P�c焾T_l��V_ޚ�t��h���ڸ������)�z�I ��<�c�^�F9�M� ^���itĀ�lU"�[����(�)~�G�����������~���G������gO=��X�c��d�'!KFG u��\*,��ߊ��m����x���U	Xxe���Wθ}�Cs�ԙ�"5a����o��KY=*$4$$�2qc����<%�kX�D��x�l�b�C �j9�.��mG��W1����`(r!��H��\��sY��D�ީ�{�&~�p�C7T���t�@�hL�#�W��:0��}�%u(}�8�E˃����`�$��b��"D=�X���w�1�{F)�����p�ߖ���vMCR����7�y�V�T�,fx��	@dK��t_�F,�V�a.Q�;a�5%+�S_�#GO��� :R�H��n\�{X�W��ބ�֊���^�}計PK$�S`��ԑ!!A���m����W(��%����V��N����^m�
81���/3#��U��6\Л��2Ϲ�1��3}B����'�����O�	?��)�ʆڌ�B��wq���&�+z�u7#J�+�p${�ш����(C�pH�ܓ������-��*O6U�~�A��g�Tj,�!Tk\��"�"j-X~�����Y�a�;�5<��r�����\���(�H"��W?�o��_q��� i8^�Bަ}���]	#�����47�U=��ǚR{L^C۠Z���@��Ti0����!�~P0h1)mȻ�L���
�d��p� Fg�Д��v���<�N�! �ͯ�)�DC5P����d��e%k��#�ł�>�����ɸ�����y����I�l8�����}�H���M���_  ?��w������_�2dM �� (@ʄ~���-�����`t��<MiSU��'�PXX�]Vt2A�ڻ��F�� �����w)gפa�/��"���g"rr�C* vt?6H�l0b�l���)�����vǠ+��h����  ���4 �t�`�w���&(+���,�s@ᑷzȵe�@J���d�Nv�Ӭ#�9��U�w/2��>�X@D�A܊�&�?��h��X�o�BPX9�v��QeK3h��tO�� ��!`<��$�G�CK�I�q�3�2o�Hs�di�7��K�ziC��D<R2q+OOvPb�2=X���@Nb6���?~)/���PwxI�0R�W����S�dr_�s�����!	����K�Ag:��s�"��$���v?���������3������������Z+���S@S�S������`J�|1�wI9�6�қ�Ԗ�>k͏���@}�k�s�S^X�ȫ���b�ďvۍЕj�����lͱj���_�͝��g$$����O�B��n�kQ;�u�n_��݆�LQԶO��(g�}l(D>�r�6_�S�	k��o�C4�9��������ў�=�����Y��1j��ľ���$�>�����ZO����Vpd�{���F �2o��b�е{m��+Z;�믯 �?=��aŵf    IDAT?��ׯ�P\/h�*	|���ۓ�&G%)��iST	9gC?#�7Ҭ*#�����/��'Y������3�b?�;�m޽�sɏ�� �7��ƟCn�fÕ�
���a�@eA BH���z���G��g
���K��SJ!l���v��e�,-uB'�H=ڴ����7b@�`{tzX�����s��������ߌ(�!�1�?����o,Z27 ��9���Cǿ4�����~Y����Z�> !o�6)�I.R� �(�SS9��FS3L2�^aez��&h��0x^^�s�I��G�&ꅓ�j�ψ7Bb���<��>��@=s4|��(*�98ϭ��/k!�+����Xӓ>�#^�w��<��չU�j�8��j�s������xI�����O?�� ��[|�����7�# ��ik��߉�� �ߣi����@�;�x��s%~t�H����c��+ P"l��w���@�^�� ^�W�Uu�^������@ �8�t��}���7c�ݰ��@+��r�^F��ԅ���Z]X� T-��r�)�%�c���'�v$�vbHNe�$Q�.X��a��YY���<�8��ͬ��UnS�U���p�	Ȋ��c\�h�������`�@����1�f�����v��� e|��{���O�����+>]/�D @����r�`x���Q�n�x<=/%W=����O<�#s�',[;��-k-����5�? ��3ֶ�7�ҷ	.�����_ф&��:C��YLFCf2r	�fu�D������ßH�C�E���a���3��d2%E�0k4�P9�:��7�Q��iU�;��x�ǧ������"�	����Qbwި+�?�K�:vM�\N�R1�T�IHEܿy��9z����8ǳG`qe�G�9	˂�;��7���|cS8u.c�s?�'֯�=&�L�o U���ad���������u����Q��])[Y�Ґ�D��w�P������C ����ˆ��'�Λ9�s��?�g��|���JF{�#��nС9랎&*�rd�X�&�ʊ���5��5�mH�e�A>�[���`X�˟v�Ł𔇰;���Z6$f�0���	�d�^���='%t�9Y" �!ok$ޙ�	���i"Vv���H�0<s�LW��4�[�v�:�S�﯎�d}c���	 l鷵�mL� �ѓ��8?�p��w!�f(�FN̟ߜ�8Ё�a�F�f�wo��A����#mf�j��
��	a?:�02]�U����B�?��;\?7�����M��}�n�6��T	�@�cs\�A�GH�N�+�E��]�6^�u�GD�.�ә��I������sB)�3�F:�����"H�:P���ѵ�~��������1^2���?�f����T2��vbӯ""V+�'�Y�e��Qt�u�G)�O��Y&bc�� .��2�/����\eֹ�-_CD�2L�Hh��m�1o��;m��ВXO�^�u�$�GZQ�	W�����>M' 0��/c}6Q��j^za��]��]]��GB��}�O�o3�?5G�$gC<�����\�4�}�.��u�#1OY*�Q^h�!E]x����c���T��#����wT�K��*1��������� D��Ͽ�	���//�H`���+^>�jf��0�x���q�l��h��s� �̣S�ͳE)�Sg'���B'vg#D\��ǡ�n���G7��m�`θ�"#�s�y�^��J�C�!��~`�Bw1���B �c������9wz�A(8V�."�2�ѵ���u�S(��A5�r>;��Z�C~���y4��t��֪i�h��p���^O2侁c(��c��x'+�lp�&_�n���_�k9m d�o���߿��w��>���������8��y{��펴'Q�(f2!.����Ï�<EE�c0�!�܋��jj��:��+C���I��A��;�>�n
�..y�>��n)6�2�d��8jGu�"[��nQ|b�-���b���8��{��PM�|����'�皚 �k���%B6G!A{��pIU]����ڈRslVǡ��պ���}I�s�_�)�ń��=��p��t2����Ѱ� ��S�j��}ξ�D L����8���}<��q(4�{RkR�q/�5S�8��D�9�ҍ�g����OT�(}ql0���יd*���/7�){��~� nS�L�ddԒ�����bL��6(�mzY�z �=��m����U������� �csu��[��km`��@GQF)���\���� (�#'�c>�3�/c�8 �}��ŧϨ�kF}�������Ok-�>��V=?'Ԯ��M��d�˛��L��G!�)��0~?����e��3�FD
���N�(�X�(0�p~ҴaK�\�;���f"���#`*&+��~VTG<��a`4[�C����A�$���]�l4�Y�.Ӧ�� �/D�5x��3��M_�Mb7�|�a+�\2�M�Z3aۮ�ow|���?���O������؏#BҰ7�&��Db��j)��Г��:V���Ε��2��o�7����T� sz|�ѯ
r�z3�	������d�O)����T�0�g ���p�W��M�A�����Ʉ!rNȧ�4��1��V Uq;*:)�:h����kD^�;�q[�m�w�v\���-�{e�&)��{1��[��rG+Ӛ�Z���7A�uH�o � ��#!���<�&�,0���4��{/a��Ѭ'p�s�&g�Cာ�:V�8����,_� �FN"c� G�q��6J�z�f$5�F![���@r�ndC��)�3��r��'�C�^ �q��������C�s.����2��p�j!������m~���UeJ	ʕ�v(�a�	��
p}��d'EҎ��@�ݐ��F�M���^_o(e�W�A T�+	kp� �2E��e�N/�~p}̏9釶QU2����5��y��uqxӣ9��6���l$�f� ǫ3�u:h�S�CDS����C��5��FEŪ��<�Wk�ð�X�xU�R�c�h�3�4�%��P�eq��r�U��9#e�`Ab���H�C*%�����C��gh~�ךnI�y�<�4�i��B�?��ӦV�D���ؔNY�x ��<_��2B�u��@Ҍdeȩ��x{�hU��D*����8�;~���Up�~�Ӗq�o�����M*����(�-���o�7q����͔)����n��"���
�X�11X��N�
c~�������>�IR
i���5���9��{5��L�#��ַ�4�,/_Jq]�3<
Z��^o��_��w�p����>���0�RJހ��߿�nb��sJ)�s��~�H��� ��^���A%"��kx�4��{����6s��,�� *`*��!�N�	ā�8Ѓѣ�M��`�9j��<���T��x���yԿR�s�<r�u�l���b�9t���@ɗ1oo&�a��5G��8��7t��6�@H���Z�8�;@��1��G[�E�+4HW1O�3��-����U:��|�p�^q�\����+�v��������I ���ڠ��~�7NhM����}��Q��/?���H?�'P&������O��K�P����DH�].�f?��'�Sc��*`F\1�O/W��gn�]�|}>�@�	�����I��RBEŖ3�;�U�`����0��[D�2��pH��X)j���BS�㜼K�L���ؤ�׵��]��uM����:�u�S��q� �ɷ��|r�Wa+ۏ'<����%�Q��$/��t2^�f��X��G��:���p�B�
DV.j�cx��0�^U�i��7S#�)H�\��7��c�\ѻ��^Q�	5(��\ʎ�������oH���� J�Y0�1�vk��Q��n��n��ܯ�f�J��F�HD��+U K}�\>Aߌo�֜�1ٰA��j�c�(��O��/� �Z�?B�oVӈ�H�R�V��n
yܑсDض��Z�e�L'�h�v�I�m"��zE��__��@�W�$�j}��t�#�-cC�Z�Ur� �b������y0�"�O� �Ia�����m12%t6� ��!����_�m�	�|��0i�V'�?_���.���'&��z��.��JN�k�� *�U;�E�j}�sq�C;����7���:��{+[��9 ����� <8!w4w&��$`YA Oys�'��z$�F1|k&�wHD�d�4�5���~���Q����-��*�Rr.���P
E�v��P�;�7�	��ʄZ+69N�;��b�t��Q�R
��.})�85H�.��?0~�����������"߾�A4�肿���4�{EO�����VA8�+��]�
DE[���<�*�p�s��x{1�f������@)l�A.�׾����@�B8���8'���M�	[�x;�~��M��!�ĥ�;��Z##Z�_/��}B��B��_��RxFYL�(��V j�G�t�+>�ӆD��vT��ز!��5 YpPҔ�^9G�O_7�"��ȱ����e\��h����$����z@j�&�vy�F�� 6f$ڰﶇ����D�����C___�Jq���6�����$�t4�R�ki�&Q̌-���Q�l�T�~ʢ��Z�j��:(W������|�~W\sB����\�)�㸽�W�����SF���7Ho�nL��ʅp}���v���kFM�nN$Q�lح�6����Br%�.#�'�3D	��rj��J���(g�ڑd�3���/�L$/e[rQ"�R��94-��bqmv�����jG����=�@S>1!%#�Y��}g���ȵ~��:G�����td�[#S%��ꍈ��Y��3T}���<Z�[a����g��c�I�
u%1D�n m2���D�
���;N��G����(cn���ye�˶�5#�@X��`�&��<�E� X�II�];�-rȄ�^�g���֦=�l|;1���X���`����{Mzԡ�4�f����3�@HN 5��������5�F}*���1H��V�<�bvg�9&�7�$$�<�/��%�4DҭS\t=l(ܩrIM�֯��SZ�ZjV�n���ێ������-������>}~���Պ�^���	(t�U �,��}��+/WV�\�VEp|�N��2�8�����5
��/_�HKz.�iD�fV��蔆#9RgK�%�[)���ڼn�Ѡ�[AVkt�5��>�V��5kۛ�۾h�ι�4S�L�,�h S��X�X��yڤw���!�����~�`��U#$�v3h��^B�n���;��jא����ur��}�A	V�O�����>)�T��dA�*���qR%��Ο�I*K)vл����+H�ʎe�+�-�������x}����^œ2����;Y6�#v�7�s�w�xP�X���m%�w�S���m?��%�V�/_�*LL��*�9;dvv�2D�7��:����xee����oի��$�hiN���Gvc;0�pB����zt�i'wMH��C@�Qa�R6�b���h0v���R�}W�z��ێ�!���@l�uB+%�䄐�&W`�Q'<i@' -�pOd�����L����a����Eg�5�<t�NƟ�����Q�Q�Jr)gC�W�	�w��R�ɊWژ��B�r)�̙���@C�2�q_kd��nM��*�Y1������X��@��C�L�h���-'�%#_����.mD�v��/��E-t̩�Nv��W<u����io�n"(N||"A�&'�Fo����9ä�k)��� r�#�����]a\,�����A"��+��u�:�����'Hk�>��ޭ�H�qF�*4�_Xq*�#������0���!��:��P��	�;�W��i�&{��Џ�:~?���9�v`���[��w�_xC+�C֣]�!εi��ʐ����*��_�Q�����no��!BhG�nhج���X�e���:�+����b�*wt+!��t+�NG;^O�a�G�Ct���>85$���i_��=�h��%Oi�#��-���?S��u�]����K9��^�s�3��R�ؐ�H��g7;$�[E�����=�����?����������ׂJ�g@��|ɞ�'���YZ�U���@W��>ٻ���Ul_uEw}.Ɉ���l6稛�T��:���Dg��׺�� 4^Y��jC!5ң������N��P1a����0/%$��������֎�l�甠�(0򥰋�X~	�`d�6�* ��n���_���UJ�dRS�{�n�2c�2r�Q�0�m"unPr! V���&�oZ�mh�Qg�֎InB5���`i?|���t�#�S��=x���Cӳ8e,"UE�<��x����ɛ58�޻"zjdb��m�S��ݥ�GI�u'�!g�*f^M}9���Of��o����|ٰ].��W�{�qO�.IƬb�q��d�X��3Ns|��{V
1"�|��q�W�#�kg��,m�hT2s���Q����r�GD�H�粒��[%{���mlR2��wK�Ql]$QsZ'��	*����.9=����^�<�#}4���P�ɮ/��
�Q
Wk=���V�>�?��ũ"��������+R���ЎN��OW_�L
�
��=w�����m�m
	�;�c�H�YF��wr��⬐W�;Hڜe�а��L	[[���������t�9�lK`�?���Ѕh���'B�l6�$-D_��$!� wq�$��pКF�ŝFf �j��j�E����Rz@���NJ�/���tD�t�_4��B��gFm�VP��=9�UP;Pk�M��kԓ�uƗ�}�����?~����p}��=���"6~� �����%!ӆ�������_��+Ralϟ�~��k��59��q)c+��;v��y���~�z��@�>�G�A:�<G�	ˢ|�Xc���G]<%6Mq�!'����>���x�c�{�j�20[�[���)[��!Q���& �p޸�U����Z|'�ӴI�,(%��C����T���n�òH���%  �¦�6'���vTS���.tS1������tl0�8�h��~0�G��ē�~�	�l��s�.���n2�MƲ�b���4Xsw@�O�r���p������`�B��#��tf�a�TU�����C/ <�[�b-.�*���������cs�`v�}���}�֛�k	�(Pjf�mD���H��QG��A��P�H��&rR������U���:"^{�1_7pD�0o�G�?F�M'��b�/�#"Pɰ�C�L�{vܳ�l�M���KWψ;��#Yo�X��&>t4]�?#�A:��%�X�~ԄR.#z#��0N�d����
��i��"�D� �7�'�!"U�3�S �
��rV�^ ��	��=�T4D����{Jfs_�h��4	�W��M�����e�N!�4A����tM(�e�٧���a�2�w���Q["�۽/��X@t�S`����v�5d��;���\	�}%Tj��u��%� V����S��s��R=���t�=�{GZ�$|w-�ׯ������u�������G��������5{I�m���`�	�M�	9[�����/���ϟL`��$ŻK�gs<,MN�z��A[����L~~�th���=��e� �X܃��8��qI���v�B���M����КX{�����g�(϶`/��`�QMHLE1S�38w?��o��[�G���¸n	�-��-Q�+��|�ã�Y�b JJ['�~1T��M~J�����(*�>�4Q�l W�ƈ]�������<�D�����H,~�@�����q1� H���1���@OV��<��LАMUjkh2�L�+�}��W�8yJ#j��K���'���eÿ�"�c�H+���Hv�����E��wD� �!0�-N(T����Q���tk(��(g|�� �͌��9D@�G�    IDAT����q�;%1T�WTj@�Z�y���Z���ώ��$M��~��p���֞�*�_���Y������ޛ�o��*�0f� 	RA�� �35Xnw˭������#��n�����%Q��E�4e�@ A��\�B�oμ���?�so���DTTፙ'��g��Z����%d�����f���++E�<��@���e��ΙJ�N	��x�(�-����H��b��(�D<�"�C11���si"����$o���=�U�7��RbYK�w(�l��#�8Ė��ere��5�������-I1Ns�=��qU�F!�7�Ij�#뙒/���_I���z����~Q�Ȯ���g�����9G׉ki][����k������X��F8:C��.��|�b�$v���j��ҩS�Nˌ� ��)$NNjC��W�`�4�oٔ���� @*3��d�Jb	�Q0�E��Ya��=��񐉃��TN���IeB�O�d��M��y�%�%7O����xsE?|�U)�^�_��,D{���Ɛ����9�@/���\x!f)�r.��cL�Q�s2k{�'��G��k�`�}d�{Z���*���I䌳���j7���*��J,		J��i%L�`�H��2/�D�c��Rb�9I%����5���MJy�k��R.mY��Y	���ȧ��Ju@?V�h���@�$�2�aб�7A?eY�5��M9c�*ci˔+�����]	��\���e�ð�Fȕ:er�D%)��W��"�*r����5r�����VT���v%Q\MІ�D9��=���4�H���"Hv�u�ʾ�=!�T�2d�ҧA�h�p�4gxV���uA��_�V��yK]�����]��}+Iu�H����L-���șZ��-���?�\����+}�qK#�
�Q����	��(W���Ң�����,�򸏼/�v�fRa�jm�@���.�&���Ƣ�Њd��^���*M��d�T�2�����o\���9$��A��9�2vs��n�.�T�ͪ�x(�w�c�Ab(D�jo��@���S�^�w�������[�G�z�cK��j��"��ȹ��=��f
��fA�Ȟ�GT�9b�xϨ$�&i�*���e,m?[#�ؗ�01���<<T�x��H9�"g#�v�$��ϱS���:���]���b�jl������Ry��AQF�u��q�6�Ƅ��A�N�\�
U��9��9�����!E]�I0�ދ������:�q����~z����S	�Y���Z�Q#��Qi%z�<f�r�+k�V�Au��� ����!����s8�	�b�z�P��q��L,��X-=�a����(pD�5o��U	j�3��a_]�d2�J%����`(�F�e�voP��#X����u7��q�k�[>��ɱ�~���Ҕ�RnF]d�F��L��i �!���ɒs�hg%����s$dI�T��	��^�	��ԋ#b�!�:Qa(�$�i�ƩY�@6KxsHb��I&,�e�� J�D�ܽ��)��\R�$=��8�E�{�x�4���;�Y&BZe���,�W�+Axx���P�$ic��)1F�V����YUܳ"k�Eo�AO�@[*��NK�_E�R��ɑ�[c.ܙA�b��K�	�f6�-}顂���Ј�Tͱ׿���8$��JK7%���;���K^Id(m�j|�$����-4a��&hBIb2g�*��p����9���P1��ҚL)��K�*��.B҈��P�etц��a!$ű��h]�,�H��jxoƌ� �f8�Y���D�0F\=��#�	�):��R�"q�j��S�mK��
AȆ�TP8(r.�EjJ�"NY�
eN��c!�j��	~Qΐ�:[.�}���LLU҆0)(]Kԑz}����=*����ȽQ���r)Y��'��Ѱ6�h;M�R�*m�1qx8'z���W�,�S�|B�٣�������6_n�(w�$��J~�[��%2|o�I�p	�T��b ��
�Y�3B.+a �iip��@����R��D�F��-~ޞ\�'uU	�Bi�����1ȥTY��m�p�	^�i�{S�)���)�l�M5��F�y�QG�jhdH{����\�:\d�(����*"Y��TW��qEv��Y�9f��r,y%��a�[Y���Ѓ-`�@�I���<��d�+�����SGf
�F���/�䘢����*�3YI`WrX2k硣q�h�c¤�5�"���F%�DiP�#1&��*�i��d�)��,?g��VL���@z)�d��>�ՊE�cQ��`�Nk��ֲ�]𘪆����S�!'|�0N�![Ȇ6w����P�PAz���$����"�6���>�HtN���7�*J^��A������I3S5��a����(dWg,:+RL8���E��⍭ѵ�hs��iTJ�{�F��T�(�&��GbH�TV䏊�"U!�TAI`����%{�<u�D�Ӓ�1٠�.L� ɷI(-��dxN
��8Q9�xmK�>}^��S��N���P�8^�a�&'�DL��G�����l�o��]���YK;�IJ���2��g�$�iI�M��K�ܡHڢ��ԩ��J��1N�m��3���1�
K�%�I.zce�b,4mI��� �t�R�B
���LLF����Z�X;Gi�h-}���&��YE-S�]*Ð�i���Z&I^w�jAnb�,�sы'd��jLt��F�@� �۞*��e���wDև��PV��i�O���p�{�����n:u�X\����*1�-��a�yْp�A��C6�d5�]P���Y�!֐z! V��$����j�pDB�+{�8��1�l��8�Q�'@I���"y�r����m��b�=,����>����I5��E�Xs��a��.=��Ά��@!j���JĤ�}�-Cob)tU����dg���稲0���jP�%�e�����-�2��3�ɥ�Υ�Py�ͬ����죫�[�j��1Xw8�P*���J
��2�	}��UHYL���Z6g�^�g�$0�a��rAyO�����laŖD"��i��c���Tr��i�l�D��(����eA?t�Ţ��f|�F�XG�V*cH	B��s5�L��zR��
)�i�5���/<'6Nsxx�I�3��[*�)�&*m0��͑�"n�r�[�q��:E�z&MC�,��9B�1g��:қ:�BB{�tNdjWs"F���]���|$j�:F�2$�`+A<���곐��PY3�,3]Ѧ��T ZS7		�Yn.Z�U`ZA�ʲ�=�d�,	����.���zzd��*[��%`��G�s���ڢ���~��΂�D	JF+�0Q���Y����@Ohm�j*�6��(}ie��i���b{�3��6�U��eV9�L�C��Jҥ��Ŵ.���S��H�K���(_�A"8�2o��@��\QJߎ�V��-��8&�S;�w�0�]Ɵ1)=g
�\��L�Lf��q�G�:]8��AR�=�d#�<�Y�|L!�*�l��<�c�fA�ք�`6�uA8�b�QH2s�T�B�D1�q�,S�Xt��	�(e͍�;(�9uz��j��gZUԕe_�24%�1��֎�������L�
�,9Gv��\����N��~����D5$ʜ(�d�pJbf1�	Q��i�i�tpi-��g��mm.NhÛ;�"n����Z�����2�L�#��K/0�ю{94�en���J�*�_��0�� ��e�Gq�*>�0e����q��RY�N�@IIHXՑ�K�?+m*re	!� +ĭ#�2(WC�K�~��]������,�{��}��<�6o=��9X��+!��oXl�s�%[!�iB�mЌ�G'�����E.'=*����,�n|=ZK�u�u�A��L�+?hx}
�Q$���H��{b��P���_�"�]B�	>���)��)b襟����zʹ��!�$]��	�j�޵���&��^ ��`�Hw�SO�D��-�G*�p(*}e��4_�%$	:�����F�$�:c+�.Ěd�B�] $/h�#mچ.J�`G,]�醘h��m',줒�+A�Z��iO� ��s�O�]��AA�b��!�H���vt}�s#��g;��C,գHR�2����++����*T��l7Ɗ�%
��\��Qs�} ��YN�q���%�q�I�=�I�ƪ��\���0��pPC���3�u&e)8bX��r+���F��}����l5�S��Zk��۟����@��E��2,�5�^�]fpO9���K�@����27^~�� %�TB+�yzx��:��g�Ť�R� �t\������l�rZ�QZ�2�:ĕ�^�:�U����E=|L^�Z)��6��隐"��SUM�ɩB���`Q8�kWn�S��֌��M��}B��f5:Ɉiqf4�3h��*�,8�ޓ�e�c��F-��fss"�LJ�$i��s��"�T(9kr�1�L�h����#�5˻euM(�(�\\y����hc��F�����pІ9K*Fbg+A_zE:�q�)�)��*��ˍ:�ڇ�/��\�]߳�C2!,���7	�d�N]i��8/����k�4Ρ�!$�<��~�=6z�F\���@r&�Rqr�辕+���@�&g�@��-a&Y��v���PW�`U򨦙�m�&�	J[�N��u5���G�gmdʞ���x�)
�8�1��8G��E�&ɖx&�uuU��y�K�Qz�37�$˚�(������MQ�eIHjm���!3�s��O�IE���8��>���
׈�ݼ�HYa�
���)��g��(e����꘭M�bb>?B�$�A�̰�õ���p�[�"���>2k6�8�ӊ.{b�Ljl/���
�=�H2���<Ejנ�@�*�a��{�ʠtE��[�4��0&|��$���h�9�(�X�HJ$)VF��h����'����u��*�!2	GC�BP�.F��ւ�h$8�{��:�2KR���".��T"r)h��8�����^z��J���D�0�E�Q�)J�L����yKNYZC��a�,�>�9��z�qHj����Y�>�c�+c1	���Z�@&EAܪ��>T�G�$n�Xi�(%��z��X�q��=�]�R"9�+D�,kd�Y��'���^���T���
�V>�!�&1Y����h1�,���-c\&�޲��h���%�T�#��"K�m�c�X'�R��t�.Vq�x��j���<�Q�T��9&���2kJR�9J��g*�y��+7�����&}��`~�lcJ���:EP�Ȝ�EY[�7�T�g�h�}�R���"\��O�l�LfT�r��O�=�3e�\�H�b/?H�T��iuݤ�A�� 'Q�x�9S�c*6��)�.�2Xu_+�x�d4o~Ĕ�!���V.��ʳ�PYq�S��?0����Hde�Y���ۀ��&���<�,��Jklm�j[�+,�e*�Tj�fJ�����yϢM�w���t*�Y�X�_�����WMntF�6G��
��0��м2��u�47��]�z�i�(��dڊ��4MK�~|���+,ڀs	�K\Q��sɑ�GR��.3�&�1���!�Z)*�n��D$I�Q��LT��2M�N,6��&0��'�&'��-1���`�[V���f2�d��1��
U�:��ts�ߜ�K�k��4�&��o[��'�ln�I+�T��vi��Y�ƹ[n�M����۞M�Z��	&�)&f�B4}�$����Cb3���GsrJl�X��Pƞ�v���uE�p��������N�>��.Y�%��r�jp�Js�=�4���~A���k���o�`'uaF;�^��ڊi�������dĩ��={�P�ơkCT�Eb`��:�D!��"_j����"tR%ZC"�A�B�Vӻ
��,�!0�I?#�L���Ge�I�k�@1ʢ��1Y��q��E��9�3��H��� �-Ҧ��9[TR��_ι$�r㌭	[W(BNYZ~9/��>-��K��%28�D�q�������~ �^v:v�k`���v��~�����|�mE�̊N��CI�
�W�i�]����T�I'ȕ\�c�8ĶRh2�^٠$ ���-�՜W�F%�ə���Ue�T5ދ߂Q����S'�qLfR|KH�J�]�l2�Ϟk�n`9���غb�pe�g�3��5��й�jI�
��ZGD�Л�lolP[��jFjgI�F�CAŴ�2 ��f�` q�{5�Y����a�/̅ݧe���f���^L�fơ!��m�̌�F�c ���
�O�@��N�9K
Yz`9���"Ӷ��7��#�J8�d�����ZAAHe-:[��/z�">$���)�g��Cb~�`~�-3�Ĩ2�h�`�mJ�RU'bX�W�	SPK2��V�ח�B��.��a΄4@w+��4���"��9�e�1��q���� �#C��V��B�Qe�]�n�r �Pt���4���=�k$E_�u��-�QPk��8eXsR���#��*Ƅ3�T��ӷ���Eߓ+K3m�)�|`�5��@<�Ռ���˾���`v�,=���K8���2�uSr�Z���a�AEΎ�F�ͫ���mS3�pp���)�ٔ8kH���&��h�F������H4��ֈ�Ȯ��ɔ�Ye&�|A�.Xs���k��ޠ�7�.�X�i���t6����� k]�`�6'k��U���d���6�����T�#���!����2�\�$#�`�W����1���!K�=�=g�ħ��Z3�08SIB%!���ʚ�����V�W����,�������κh�k!4� -��\(%��2�e������J��#h�I�=vR肶h���x�}�Z���4gq΃"5-��#){���!���P1+��vz99r��1J�g�j����Z򕆷�V2!T�Y�V+���"UČ��`BAw�R��r��I�8H����0@�C[v�������)��%�:�qU���c�dF��>D���\�T�_����X�+��k5m9��դ���h���՛��Y�7O�+C7�IeN!,A)��%��۴�8c9�<]{H����h{n�=�MŤ24�	��	��䈮�"��T!,k�ǹ0yl�jr�; �c���氲A�a(�/#�S���7k+e�5)�6H����]yon��j���B�JJ,C�
6C�˨ٶ̈́\�t(AJE��"��$(e�>�"�(},�DTRx�Yt��6���0���R
8%�R��Qo��W�J�ó
y��i���������.���1�*�M��J��p��{��-3@熬/@F��c����i�<W5؏&9H����#���l�=��?9k���9JGX��(�G�>[�֠�����G�
j�YK0��.�z�b���v!6�1���ٴ������{4�[�z�N+���8�^���-���l��³3�x��>ŝ�}/�j�?��=�].��I�y��;`������_��C�R7kh���e^����������r�ּ��1����n9C{x���'�˫�>�y������d����9GJ'�}�	��^fۛ��\�e^��wY\��&�^��[�������3?�}�"�e�y�[Ǿ��b�>���s?��9�k\z�2��/���+ldM�u��!Lj���Fۊ:�)�aV�a�9ʙX9���!01�Y-R�6��8��wc��s�iÚ�h����<F;��x4��HCơ�*�v��*c�C ��9�L�5"+~�.��Q=���\N�1@֠E�)�����*-U@�TV��{d���5��E�ŭ."oeRA7��A�E�Ҕ���H��z���C}1�)2�Q���k�IA�2z5���n�_>Hㄸ�����e%hj�Ę*J�+�����K'���g
O*%�72�+�*!,EN��5�_��"Y__�6�)I�UZ�H�mo~�o�f~����M��&',�5!fQ|�J�Zi�ʒQt����Y����/_c��&ӵMZ��HE�,��jhk+�3ð�^fH��/"��ɳ�Ym%q��!��50ʎ�$Q�?�"rH"����l�x�%F�����7�m*,�qqWu���|�2�1�Vn@[p�z��     IDATଘ���6���{��,�e�=�6�{�65Y��ٖ�hT�n,��ᜥ+��R�rN�8�e4�4}�8j{��21�~����we�i,�T$���ҫ�Ky�ƌ�;s����� k��ZO�b��G��<^��v�T�*�!��Fӕʊ���^���a��禜�aQ����X2�㩉*WB�D�JKBB�(��S_*��r1�����d��*˦��c��c?f�j����O|�殻�M�;�0W�s�k�`���qz}5���&���N�Wg��2��4n���<�7�^C���9s����>��'���W^�|�W_��~]��눽�N�����U��6:+v/\�c��~v�{������=�m�?�#_��>�~�����H���~��������+׸�����4�|�#����������������(g��S�ж-n{�{{w}�K���,vsFUk��>?��,O�ٟr�W9m[g���/�����ޜ�^|���Xw{)b��<��'�����ؓg�?�c�������^z��[O}�$k��f��yt�p�S�l��������O��ݣr?i��&�m�.^�?��ێv�9�Ʈ�ѬO9T���5��e~pH����11IU����Ja�60V$Q9x��z*�;G�#� .@ѿI�`��$cTS[kce�h��H� �G�5�D�^�Q��Zx}���(*�&E��Xt=��(�H�2�������n�s$����Ȥ�@ʕ�J'r�a)���=���ἧ�8h��o���'���+�ᒔ��3�Wk��d�(�;�{�E��Ȝ���^x�\~W��*ÀR����Qf9gp4�1�����V7�,��XGU�+j�Tc�0@g9b�Th���ؘM�8}�����>)D�6��z1l2���S��̦5��c��7�a����Ţ���[�>q���ڣ#j%fl¼T�h%{�6O�
m�iC�2k@"����*W4��T�2��D�o���8��	�X�/?�J[ehK{��� �:fB��WK�WIzLZ)��M�/(r��Z�Ԯ�{����D'��/�TMS�5�2��d�]��ؑTBP����|�w��@;Hi��n}�S;�lRaj��d�І�BU�X�-��`����Q+z|�$�I�}�6f�x��C�*2i49�K��У*ɏN�)�h٥�&0I�*r�%�q�
#~��Qe��1z�e���c�R�v���J�P!D��$��8�bMqk*�G)��y��	��r؄F�d�+O��:ҕ��=�T�z��ҵl��<�?����9C�����)w<}�y���?`著�=���ſ����iU�w7�ؚ�#�����C����k���O��~�jcK�*>�x������������ g�|���w��S����O�N�վa��q���n�s��ѳ-~���py��� r��f�>�={�Ǿ�.��qt�=�y6��(�_z���_�ԩӬ����x��z�������OXo���ɩ#LZҽ��¯�/�q�n^e~�2}��4���A�7�����W��'>��<��������Ѥ.�hNq�]��;>�[�Zw�������y�_�ǿ���N��_彏}�����y�V�t:E��>�������Wh����r?�����<�/��7|���-�{�����0rE5���/���/鋸8a�n�Y�ܳ�����X{�
�eK�m��5�}❟�,���J��0ϥ�7���7�ug�Nk�p�{>��O?�l}�~����n��3^���p��9�j~|��>���YO~�����f��R@�6W�6���ȭ��g�&;��v�v�e��_c�{�E7[�z��S��q��â_���S?��]�o4\ٿ��n���G؊��kv�`��s��	B?e�G�g��� Ѩb�]n�	#�]K� f`��@�z0^�Is�{"#v�>9g|7k���W/ڷ!���ּYY%?/��"-�֍AlEʚ.dj�i4F��I���p�e8$19ʰ���bņ{�*�l���AZH�)Z�|��f���>���6�����1�
3]��KR��"F�Ɂ�Z��.��ZZ�֠7�� �Slo���ឨz�H����Z̼�{�5L�
���ӶN�>F;�89mF�$@G�*f�J�Z;����9Cb!"k��Q+q\�$���)����E���2K��X͗�������x��j�suɲJO����h�V��t�3Z��L���	1ѵ��zOR1c��9�VL��I�+-��x)��Ӣ'���6�M�|H�)rW�����B<Js�5�d��r8V�������B&FGJp$��稵f�eX�l�$,�T����׏�@1)	iU�ddE��qP7�J��]���������������ս�٘������w�/�:�.�ŋ�=�ͯ��3��wr��>��m��K�'w?�0w��Q�þ���J�:Au�=l�y������p�:�m����������ₓ'α}��}�q��_���\{���ml�{isµ~�S��|�96���}�]���&��2v���ғ�������?¶��W<���	�}�W`�ŝ�?���.w}���r�"������g�C�?���;�#Ln=���6�JI�}"�}�<���7��?������E�����[��?�x�������Oos���hgIܹf�yl�y�'T���w}��4�-���п�
a_��������'>ƅ�a�%z��l�;�����]~��8����4O|��|��_������<���Μ�p���)j�BŊ�l���>�c_�5�ٜ�'o��	{�-��<�;{�f�x�������T�浝=���'��o���n�7۞~�q˹[��y�O��4�x�W~�G�k︇S[�\������2�V>��_~�x�Q��?����.q��3����(v�Z��^]f���㷹�}�&�L�3S�y��g����0���h�{��}�㗸�����{��}&���k?���O��ty������'��s�g���f��l�q����C��W��Sf��0f@�2Bz.@k�۞����/��%���z���1���!�UH�{A@sc܈((�Dm�	
�T���8���RXS�?��20h`�(����#A�Ǟ��A6��9� ,��A+�����v�9o��y���X��2�F-����9����*1�)�G�2���@�/��;w���:}���Pi�t:���t�B�N9�G�X��8:���깪"��������&T͔~�
�^+|AG\U��Od/[���#&sL,\�7u5Ɗ~x#J��f�j쭶�)F����^.�߆X���IIU%�\r��`Tq�+>�F�1�3�7�}�me�m�r	̔I�Tuʹ��+a$'�8P��d���b(6��`�1�Gay��眄)Y;f�H¬Vh#�C�����&�6���+LZ%�����2�v	�����/��(NhC�5)I߭�/룸��2h���8zd�co�� ��+�A��׼�VoV�N�5����kx��'ư��[γy��tNsp�?�����W�n�A��u����� �[l{��g���^ϓ������u�N���������lms���\{�"��/��+����9���<{/�~��������;9}���t�2'�	��	t�0�V4G;lܼJn�x��_��o}{c�I�G�������ĠiXu��[y��e.��0]K\?<��]w��Q���K/s��U�\���}���8GU�Ʊ�JYL]�]���w����^������0�
�}Y��f�/=Kz��ŝ���}�)��Y��cq�2���܅;�c��^z��=�t�]�'��X���<��ٻ�`��5��_�/}�[�Վ���s�|��oq��)n{�!rS�XAH�Um�^k��� �������y��'_�
���S6N���2��?��'~���~���78�<�<�(���/1��vvo�Ć�+���v�{~�O��?�������Я~��|�K�/b�w������!��u'���܌K���W����5���}�Ҧ����S
�>D��w��|��?�k*v~�2��4����G>�Gw�����A�j>��g��N�5�"z�>��gxn�g���'��=����6�ﻗ���#'N���S�c�ow�5��x��Β��,�Y���^
�6�Q��J�]���]��c�RǾw��cQT1_�M:"���B4�C����C��&�J�
rz%b�#ypPr)%�+�JP̡�P*R17%�q_�b�%� #n��y�k�^��[O�6���}K�rkP	�0��E�����8��4zJh��ve�|z���'QJ1�ۧ�QEq,��Xm�
��2�����c�%g��|�(��r��E߯WTK*��i�
+ne�xl$�����!}���I�h���Y�Il)%�/������/= W�����:bH��t�G�0��ã^��A�U�Rt�fb�M*�J��~@ ��b�S�~�2�lh�@�fI�"WN��Sh�65�IMe�}+H^t��C�2�?~�
�����e����,g��68j��膍8F��Z����H�3�e�Ġ�l�t��N {y��ؔO;���������0f��8H�A����m�'��8��6��1s{p�N��޸�w�Ϳ��S����%f��~�c���7������:�5�G�̻}n�	}����U^��7���bqu�L�t�)���p�/��S�'��r4.�U��Q��U5a�4�՜�4��c�s��l���6�����qb�);�S���Or��>D}j�+��/=�c��»1ʲ�>c}�!��������т��#eKek�6�.��C����mm&���@=es3p�[�7�M��`� �_|��]wS���ȡ���2��/?��g���p?�������ǆ���}�p��wC=ag� ;��6��L޻I�z��2?�^����xe����Por��1=y��SSf�O���8p���n����l���&�lϘ��8�x��~�=6���w�No;Bw@�����}�;��Nnܸ�s��?��W^c�[q���<p���u��W�ek��W~�w��G��^���L���?��y���}�[�=|�s�����U�EO��Dc�Y�miN*�.���cV+���7��_}��y`��{y��>���� ���-^}�w\�����<�wNz�u�AOw�9ο�ݜ���?�0;����?ȉS���w�/����	7x�s�x�<�^��k<������W�\3��Փ4�,��\Y/��۟ͷ;�ow鏿{%f-�D
0*�+-

(V�����M���Nȸ�]�]�0zH�Ń ��4�di?�2�	,�O^�v@�c�Ru���$��H(��s�Ir}���Mn=���t��L�%��Y��|)�,�g4j*E�|��M�lbg�s���9���	���-��RkKO�	�k���O]�Q�|�Ĭ0vJ֙�E�W�[��8:أ��X��`��T��T�V��eT�T���Շ5�(��#��6ƱgH>��>F�V���:aM6MEU[������$px(��C����,:]z5j9w=G,��f2�����������w�y���Bf>o�;Fs;Ȃr��DS[f��YUl?���.d�����[�V���N��!��?�o�Y�v�2�Ojb�8���e��Le�ϴ)J\BI҆��#gF�~�"�+����ҁj�up<��b2�6jPTȘY�*|���w�N@c];�G1ٞ��W��)��gNlspc��+�4vJ���['x�3���;�2���5�Wa�*}��Ln� 7��=����g8ur��~ʥ�_ �hei}�J�%�J�c:�������2lO�i��*�����~��[���3��G��ثװ�CE`��͏8�-���}��l�3��Z�*HZ�����P�s���^z5�����{g��/����~�Z�D	��*E��˯<�O��m�w�A>��g�:֫)zn�d�p���looR'E���3�ºs�����<C����3������!�x�cd9�T�ӧ9q�}�{�mx���/��4g��]_�"��;y��6�>�։m��_�۽�Վ�+&�T�5^�9?��W�^�9�̯��S��e~�������ȳ�ٹq��g���Ϲy����ǰ�3�6gp��E����dr�^�/�#qlt��8w�}�A�{6�i���2���?d��"�)��}N�o�s߃0��R{\z�ܸ�S.}�����P�μ���_�v�>-�jA�����}����?`q�i^�����e>\Mx��'x��x�k�uc[�/��{#��3��~��/"�cj��E�@�[��Qn���c��3F-.�*�C��e{]�N�ur���5&��������Rp���KH���\|BB��H2sbq��8ƛ!v#yS�hS���e�r�{Az�Nkn��k봋׮g�uM�:bޖL�Ћb?��؃O��-�DH�E�\͢;�׮r��&�Mt=e�&Z	�<��̙,�]��Ȋ���.II_�������u����D�2(�R�p%a��	J��7_�ח� .�hC��Z/�h��J���v�D,��q��t�1���[ ���-�m�98��z
y`�Kժvm����¦M��a�T��4��4����-9�Pi�hS��$�ڰ6�ehM쎙����&��ck3.����}�8Ō�
K���h�ٹF�(5ZM��fIZ�*���ب)�AI$��x�����5E^���ˡ�{���[���[�vx� !q��������4kL�#�[��WMH��!������g��]�3q�j�Ƒ6��x���>�9&�f����+~��L�&lmv�ܟ�7;ǝ������y?���������{�v���6�4��!�9:vl�m��ȼح��+M�n�p�'?��O|���S�7�`��|��o��M*�V��9��3QS��r�R�W���g�j,����Me"W����H�����U;6�<��3;/^�9�B�l�l����K��G�}��67*M[5�p�|�eۜ_�96��e֔äHT���b֧�����דd�y����1��u�o��	K�Z��(�Ԉ�fF�������^�^n�^�_�&&b6bcCژI�D/�I�
$Cx�э������NfU7�ܘ�MDG���N�9�3�����<d2��ң�wo��2o�Hi8u��;����a���E���q���(��y�Ǩl�7(Q�a륟"����B�O��ǻ��+eK��j]3��3��f\����k��XN*�<�G�~���1�Yר_��_���O|���s7kGNp)/�ن2+�JSAA�$�ر?����ð�Y[r��u^�OK�}�."�����Qm_d�U�R�Z�]��0�O�MTs�d�^��?�������;��'N�������S�N�*K4m�[��u*B�~Ym}�Z$�2�ņz8(8��M�^��%���ɔ}/J!�RċHT�� ��戲�̧�L��x�24}�˲,@�Sp�����`�@�N2�~�%Ow�a�hh;�����01.�<1��6��y�'2���L2�!���AD�2&%">!J�4�E�(à��ڈ.�#)I�x���Ǩu�׆��3��B��I���:)b�p!i/���Y�hmC$u%ضek{�c'��z�8{7��V3����W��m;?��:1#�A+�-M�������m�:AW�H����b��5B&("��c����)hm2��k��*��u��R$�z�ѣ��@�����:F�ka�x�5����b�e�΂H�|��BR"�$P jRݨݠ�N-'�ቹ����@�xW2�X�5D��N�)��}����=S��2!��pGt	� �_�r�ʎp�N��V� �[�����K6�_����u����~����7�M�\#K���6��͈IS3�0�"�9E��W%7&5[k=�����o�.������/��~��9GQ�X�pa��cO�������ٻr�����s��C�J�K7E�@	l�״1c�r\e���9v�}��=�7��+�UN}��|����ͣ윿�O���\}�_Ѻ������\�d�Ĭ��~�\+����ꏿG}�<*�o�)3C/S��)�%�    IDAT��Uv�}��}�ɹ���8��l�*囖#f@�*��vV�\ ��	2玻��>�U��|�4W/sdx���S���cl_��{���H]WT�);;;�֒�
jgP����
E���錙ќߺL[(��S^��yn{�z?�x��[��;X�\?��9u����a>����1B��i�����ٜ�Q>bV��"8��F��?����|��tɻ��#��>�訂gP�X=}�<�A�y�;�/_�H���r� �{��gSJS�"Զfg�K�4�8�lf�Lc�7}��R��3�#g������(�7��.~���B5e(3��~������c�\r��y�����e��J��Z����.��ͼ��'�5����T�;��ە�k�-��.�;���z<'��}����B�����}�,ce8�5-�;�E~)�ە���p�[x�,aɖ�²ĸDM�l|��+y�@�-k���ܳ�?'I�� �E�DB�LC[M����򵌝iW�F(�E�ܪZO����BPf6�l��EhA4º)��������5Pj�I
^�@Y&Ѳi�Ҷ"M5o�ٛ�2C9\EI�uU2t��im�1.;����^'h�����f	�gq���2E*>�TI_�3� ��Ki6���%F|T՜ɬaȲm;?�Qˤv����6޳�8L2IpQr��ז�������|gɈx�5�,Ɍ xK��"���V���$��'�AT�%���6T�B�39tJ�0��t��^�պd>C��4:��]�WFỚ��R�A�Y�.�Ӂ�Bt��� =qK�p���b��0������{���E;�~o�2������! +Olי�d<�r�ͷ���E�;�v�G>�;<����_2�x�7��%���_r&dȨ6���я�����g���w/�ӿ�[^���8�$�l�����{�i@�s�^��LkN|�I>������g��z��>�1>����ޑ�.^��~��^�)�j�scn�ݛ�7�����3�C^X;r����X-�E����%�s�Q ��|�W�W��;l��)F�����x������.�.�'&�5��&r�4�R[�0SLww9"r�?s|��q͍W�������V�X=�����	3g��F��B��M�d
���h��3���4�<f�&n�ǭ8.�r}%c���a4ൟ}���e����������;�k%���fG@��l0����O��O=�D�L\�Ɛ��628~����?c��ӬyŹo|�_|���{�U�Wf{3z�����Nb���nl'�ƒG����1�Nq�3��R̥C���Y`��pUdhrz�ǎ��18�ß�S���X[Y���>�[�U�;7X=����j���+o1��,�T)8���{d1�C��T:�p��"Yf�˵�vs.�n��o������`��Yܽ����]��7c�_����T�3hj��-%���A9Uk�4j��K)p~��Jv�A��o%S�(�,�Ӊ9�*�Z����u��	Q�X��d&g}m�d��6^H�Ҍ����"ǶslӢ"I,Iij�L�xv�%P:#˓��t�R�%v�bH���g\���Qs�����7mP�Ӧ���{��D���єf3KU�7�^���M�V�y�	�&�e9$�S�~\�&>����?t�<�|!���C�۷�	@�1Q|H.tZw&2��P-74�H�ؕ2&����N� �&i]�P��p�()��W��t� ��q�E�㜣u	RiI5o����j��RG�4�݌�0E�VI�2�Ā�>b[(�N�Z�O=��mZd7��1H!��u���L'}Ҹ^ԧ�k?��$;U�Ұ\��(���[W�	�hA�
'"�ZA�`f��!m�"�������@�䒬He�� ���9�7C8���e�qA�\�OZd�`��� � 6`t�!������|����|���}�3��3�����	����x�>NcV��{����_��s?dqm@5o�r@��Gx賿ý���ƅ7��_�5��=�}�S��
�+(����!�N����{����3�_����u�(4�ʇ�C������Y&9���8s�Ѱǻo�����Cx�'�O?���ɿ���;��_�p幟v�Հ�A�5j"�����1*�)�����}���w�i��g���<���r��D錓~
1��=�w��w�s���y�����_���=I��W�q�!|�d~ieŉu��#�y�)^����׮`O�e�c�p��q�/0��A�	��2[�ݺ���Y�>�R5�U>����uvϿ������;o]�诒ݤ8�ct�O��{!G�/�1����;�1~�:���h��ezҒ�	�e{"�ￗ������&����������9��g2���ML�g�d�j~���Kh2�8%�uͺR�9�j�KJ�v\
jE�#{�ǂ����i>�����������o|�k�a�6�5����0�����L^�f��Ӝ��Gat7����k�_:�	���X���l^,��˵bcs��pSV������Þ"]ORB�Ę-PĐ�ޣ� T�䬭�`-v��2�b����%F��H������@p.I#��բER���#c�]�wF:Gͮ���
GV���P�Q�A�A�֢��Zk�M�
A�[q��ʉ�GX;z���v>�(�u�	�x��$>@�`�y�U;�IE49Aj4���޾���,�J+����`C�+p
g#���z, 4dRs�����C)� /��ʹ+��L	lt��I�k�j�,6��;���5�D:EO���ypܺ�� ��H��Lm�5�E���4>t��ݐ�!`�$W9Z��:�W�6 O�"�e�Y���jh�K��*�tJ@�iz2i���,v�������]})q�Tx�P�@�=���;�n�y�o�:�1]m閶��"���"��J)l̓U�NѠk�#��`�"&��(�C�Ut�7��B
���?~�=�/}$��������
T�tw��7��3�s�SO�3����rG�('?�Iځd����'��x���	�V����\����󱏡�Ǳ�����^����<�?�kN<p[x�����Cw>�@¥�os����&�ɔW��m�p���ڧ�8}7a��\�8ݗL�|�W��#����O��z8�9�#h��ǎ#T��9{�1������S��=}�>�����3��u~�����~L�ִ�E��2/(2���[���*g����z?/�\f.��Ư���R�}��y���G���N5Z���G����=|��?��ƻ�틼�����Ü���E�S���9�so����G�z����E~�4�?�4�hح���#�'�c8��b�E.�q���Rek�j����|5�}�x��j��eǑ+s���_z�^���ǟ���1ۺ�؃�)`��1�n�8}�~�3<�=����9r�,��������?���+�'x�c����?���}�~���@�U��
� �&gV\#��,ֵ�K&�#�k�:x��5eV��k�Ռ�ǟ��s�l���N��(��n�v���o?Kq|��>��<���f�?�Ͼ�U��Ɨ�7�����8Ǖ���yUl2ۺBo2��_�"��*�=��ާǜ=��͓L޹�0������k���?~�M���9�!���D���d��Z�Cn4���|b�w�wr]���.%�}�� �:ą��b]J|��~!E�K?� ��v`�[�֦�-Q��EP:yH����ltc�9���%��K�,'��?\c��tF�g��g��β�yc\�e��@�6�q��9��+��JV%���{;�&��{�nj�0�D�H�i�,co:���8��,^G�N��[co���rz-;���nW�}������>�W�����z���q��Ԉ�;=�j�A��
�IJwBdg�(��EO m�.¬n��
�I.."XB2�)3CiR���ӻ����H�̓b�R��>N�ŀ�졵X/�kC�(y�t�̒}��/�XE.n&�F�sԺǩG�g�\��N��6�<����Ow���e�$�ɂ_�P�pHR�ts���&��޿x�&��n,"[W�g�z���{z�p߇�౧��ޏ|��n�~&P�m^��W����x���1���?���G2�s��W����c�s�c����n��w���am��4wU3~�9^��78���x�����.�?���m�i�����R��&�������or����L��eF6,A�4[W�Wށ틼���"L��a�ƩS(�ع�åg���_�*��-D&�yF1��)7�݋\���Y�n>p�(�GE�}y�aV�^�����k�Ǐ�#,>2	1/Y[[a����d����͓<�G��V�Bè'�v�M^�������'[]'��Ͻ~�{����cLWK���e���y�0�������;���I>��Ğ.x�{_�]����~��^Q�y�4�=���:G��u�2o���4�;de��l��� ���q����w�,�޸���q����ńW��	��I��o���$�J��kW�����W2|����W޼�y��}w��T�U�y����W���2�����HE�rFN���������T�>+�Gy��ft4����=��]��دq����\�t��׮0��!��u�z���E��O|
�������f���ѣȞDk���ZO�\��~�<Zn|�d�����[�����s�����69�dBB(�ܯ�:}R�1��$g:�d���@�>Y`��	]��*]>���Ε>8�N�-�T�R��1
�@��9�CȄF�ح�)I��:%!z���ŪgW��r��*����4մ����!x�j�<�H(iX� PH����΄P;2-)����,FH\�I����J�uc@���Z�#�e��-^����e��x�[��$��ѩ��zn\�d��!�:�D�7s�85��dަ������ɡ'zTd��0�̨���1�S9��e�w81y����tF�x�W��tr�s%�3Ead��7�\J,j�s�����IŬ	 f(��z�i/6�Ä�,$S�bRFZ��w����� (����f^��>b���޵�x��z6#f�c^謄#�HR�z:�e��N�u<L��ݽ��y77A���O@SL����'��{��+?et�,�Vȧ�v�����ϲ:�e��p^�'hL�r�P��r._�m(����M�2L�T�)�d/��ۥ�j�а�	ra�z�"?��/|�o(����:�'c�$!�~��p�^D1���mKP]P�PM�_��ݣ�٘K?�.��,G�6�{%��m��^C�Ǭ��l�'%r� d�^%{���ş�g�<��i��̷97m��_�����Y^ܹ���`�W�bϝc��d���˕�������:�� �o���7�ig��=^��_0�E�����>r}����+�x�l��s�ڈ��_0��u�F�o#�_�޾��NX��k��u�k��ά�V�X��$W����w��W������MDL[���"�~�����q��6����sV������|�����#k���C�kU�Rl��o�8�z�9sL����3����?�棏�lE6,y�#d~�]~���!1e���q�����s��iN>�+���	HrY���gy�~����'>�������a�'��T�:���]�����w=�w>��d�l@��Sg�i�]��~���fTt]<ݺ��r��ݺ��͹[��[������a���cZS����e��MG�f�=�O�J�]Y����-�:ޑ�&�[w�̙x`Ig?E�IZ"���M�Q��u؎�'�zz��Q�dD��Zcb'+�Mk��Μ>Ju�t�R�X* �N^��7(i��.�i�٤���8�~c����+�X3��LS��" 
1(Ba�!�@�ò�Ae=�� �A
�!URqh�����q��=J���gq�⡃^�0tǸ��\�5WU�n����O'�E�)���&�����:�ۮ�@(��yU1�-ŹE����^�\���K����t�zK�}�O�Z˼�Ts�s"�Us��O�ч� !�.zY��1�c�)!i|�ib��6�@���<��qd�S���3���/7��.�(R��A$3��HB�a]�u���HBD�{z�(n����	ᇮ&���{R��	��)�M͍w^����q~�@�̮�plu3:�k?{�K�R������`t���);�7�8������E$f��Sh����+H�Bbc����Usƻ���'k#Z!qY2�d@֖����F(D���H��EF��\��i;��4f��ULQ2�<�^�K;�\3��Lg���ڥm&��fV�DÍ��m����OPd������].�kb�έi�Ⱥ�T�K��_˰՘���+T�H*	��a�h��K��+��uLV Q��eG�W�I��{���/�fC��u��V�쌾p��l���M�܏�/T�̈YW���r��y�����e�Onp����7_bw=�~d��s˵�y&/�ȫ��&��g����>���(r�hif3���r����z���K��y�8"�yD:���MIpMp�L3_�܏�`c������#�v\~�%~������s��èKWpo�X���Q0���6��f����<��O~�_ŷ*����������O?f4k)�����@��f�X�o%�����[3`��OH�!%��=:���"|��Qu���Hi���6���@$����`4(�
��AL����*)��l�� 	<���~�.Q���ʈ!$h2r`T����c��X�r2�ڰd<o�Ca2�\����jA�����U�ˠej�^:�ʀ �iŰ4h����[��,�i���k���<��+�����ԁ%����%J�����d�%��%P�dJvm�cq��D+����˒��?���dw�ڶ�m�S��2ս���C+�ںao�؆B(>e�RRf&�ಂ;U;6$��(E�d4���*yHx��IhGDK�)����Ԋ�M��b�>��e��m��a^Y\�]�P8@�eM=Ƹ��ٽ1�Sj��}6�#ګ�6�Ó0ƈ��~r2�ŝgϐi�t��Q
k'hq`e��_GJM�8&�y�Q&G=!:.�A��c"�,zdo]L?�$�{�M� �;��ةv��E��2��p��G��LI<9hC-NX�V`��3�z���ϙ�C_���!�|��
CSh�c��'<!�0�60�P�C�ȲO�"!N���i�(%�vBe[�h�.o�����7�D�}��Ɔ��*v���$�9�+.\�L�/�cu�Dz������\�)M�W._�k�9q���յ5��c��:F�w��Yb?GJ�����LYt�S�9�6��������;��e7��u$�!u�h�V%�LȰdTƓ�^�ՄJv�v�i�)�7�{(eI)5s;#���ѻ3LkX��qq���26}�݋��SZiY�ټ�ꕋdF�8O�#�\��C��^_�w����}��+�{�!i�A�l��+VVi���Vpe"!��g��^������ѻ�d4\%jh�}��|�p}�̶����2��ów3<u��G��ؖ�n���+T��(B�h���qF�7Y?q��cD3fP%�3��Wx�՟�����#�c�|�qVB�π믾΍�z�3E����D%X�/e!�2�b���ub1�n�~��Xw�lX։�S���\K�%��!S
y�չ6;,֜���S�X顳]��JEZ�;Y����n�vM���)�\~�.Ql�c�"]*�Lc��[��J.p1սC�(�R_�F��iei�B(�u-�ln��:�1�ߣ�N�"���\��]��&>H�cV[Z�L�>��ύ���uF�a6���I��c
@D�kHL�DBe�(��-�M"tenȌ�^H�eM��Z!i���1y�w�������k[��(���e�!���=�|9X�t��'X�"Y)z���tQ\ ���2�����r�_���E���p�к@�VL�5!�12F�L��J	�"��5����Ò� ����C/������*��:�E����'�jI~�J&����RE*���c�    IDAT,����c:ܪB(�q�\@���45W.]�؉#�׷�����;�d��Q2�I^(���~:�s�d6��k��.�}�����M~qj�n��O����/ ��z����dVb�ŋ���*r�������>+�����k�*����|NN�P��	-^�1f�C��$�y�� /���؆�(���fc�7�\�!/{77h;���l��1�2��PBSh�x<���8z�=���[[����J"}dE�\ٽ��k�<ʑ�5���a��Bpm�CJ�DЕM��R���x�X�#t4L}�ۗ.�/{�	2����SE���Ļ����(�ƵM�v��I*��P;�PM
�^NP��?a�ƌA�$
��#��aqVB�y��96�)<� ׷v��szs���*ާ�i$u[S��{�ʈ�ic�����OV�(!ٛi⊡�g�X}��<hW1ߟ�6��z?E��ub:�CoЧ_j)�H�x^1�fTr��h�O����o�3�����f��jw�/,ż6O���; ���7�~����'9�����hn\f�4�ķ�����U��[�s����J����M?'A���<JAQj�<C������z�bAN)�K�`�7'���s*��A�d��m7�䮦�;ݐ_�aP��tJh"��YYY������ ;@Ŀ��yVuZ��K�c��������Nk�Vxپ>���0�!1
�lBm[�(-@| A� ���:MѴ��%4um�ٞ �F�������.�A�L^%"�V�E{{�09v�B�[eK����
��>ny���nya��+Į%��`]dk7���f�hqC�,�Z)$�H�\�u����bR��ZO�>I��d�I��B`���������~QP�i!w�%��Fw�а��xZ�X�P����Gl� "h}����tׁ��B�:�1K�I�A�X�,Q.n��׷
�"�eU]su�*��68s���^M��	!T��ʼkj�T�ƋԶ�]׫�.�{Z%����m�J������q��v��ƀ��ck�F��6XʬA�{�5C�GT-���L�X��52W̚9�h�¡T���h�SJ�R��'��	�'%5���8�Bm�f���ƾ�ݵ�֨���2�j�49nޢ�3�3�� �g��D#���g4ȹt��<�SE�h�|�<�љa<�"�cU�r���Ԯ��Z���,g�;!�)�b�H�M ���Z�ld�]�d9�%}m�'�`Xп�$�����h��xoq�3S�����e>`�J���\"C��-�������qOTk�6����YIa��uK^#�)��1�W��;f�#��R�����6�GD��MCF�T���)�l5M��V�s������5efPmƶ#sI�b�4���MYE�N׾�92ϨD�Ui������P�T�R!�E�mXk%���_�3�r)]��!��IPl�
���.%�W��.cw����ȩ2�+������׿ʕ��G�~������Z"]̥ï��5������~q�	wA'��� L��D@���%�43R��=��I�],
��8��R���I
�Y(�N�_~�*�,m��B����T�Ъs�s�!	��EDܸ�ƩM����n�W��2�TW���y��a2E�_P�>%HB�˥�[�9y�յ�=g�*]�z��j������&n��%�2C(A%�ji�*q~���	���q�)�+��X0��(�t<.��S#��X绽%��y޿�9tQ�]t:$�io:|�տ�����Љ���h� Z�%B�L�D,�D'��\��Z<,���������r�Q�;^�I�BtJz-ѻ�V`�~�3�5�jK�2�bDň��j�B�+R�Ԫ �Q
�X�J�bLǏ��WLf�Yd������AEH>�%�"
�|M�D:	���"��G�$,E�*':rL\�X����!$H��yb�d�Ϩ��=Z�M}��.p�� �MH}��%�X"��XH슮�>�dj�[(�(����5��������N�BC�D�RۍP
�$^D�Y�Χ���}�c{V��Z�u���(�a�@J��t�fqu��c�B�A���R8|փ���J���jK�f���>����1�R�MulJ3�׬F�(i��5�h�U6uB�@h[���F��9��,mh�*b���2Tۢe�*G-�k�B�G�D��
��"�F��\�D/�tIQ�Fz��޳����FG���,�*궡���M0h��i�W���L�bh%�d����'�&[m)��m@*I���t��✦�`��y�
�B�	I�޵T�/s}g�>&��2���bҐ�M���&�Zh�������Ϻ��h�3lc�Qqm��<�8穛
;����� Uƞm���N�9�����.R�9u�`�}�B�o�U���	�)�6���A�!4�U�Ԉ��IAkF��eNi�~�y��B\^b��b������sf;c֥"�kB)���32%����E�ۑ)"J���HXh��vZ�j�2=�� e��;���<K>JF�K.$"ʔ��ź�=F�>�ʠQ���	ε��"��dC�F��]c�&*��s��i��RР�B�P]v���?)P2��h�6�$&Q�ӾשlidDZK�7F��<u�w�@Y	�fE�ґ�����QA��D������PW� ��)�>8�udQ�����v�3J D �&�u$)�|R���e���`m��"�o!�lۡ�
#X��@^�~���C��2 2�V��d2*��
A=����8�k����$Vʔ�/"(ՙ�I.�����"����ڼZlL7E� BGIu�[T����B%V&
$D�t>�j,6�4p�χ��
my���!HF	]�A*E�}ڬLN 	�4���.3���([�%�u�&��`�۵����0�X*�Ԟ����|>���&+p61cM�#8Ǽ���|�#���L��Ȉp��N�Ȍ�vDb	J!p������#t%�e��a�������Npe��<A��(M�Λ�]٢V��.:�N�"X�I���5D]���5�����JCM��C6@�-r�N���S�r���&C*�H�>�/�[�x�����9�O�u��dX������s�R $�h�#a00�L0J`�<�Y�P75���H��S����15�LFM��#>�r�>���*�	�y����ֻWY�(h����>�V����z�A�Vx|��C�m�޲Q(4�j2'/��k�K�sDY^� ��7h<jZ�a)�����!D�;���1�:F�G(�ّ!�xt��H���3��Xߠ|$J��\�!��Yݰ�w���8�v��"�&����"�@?�r�LڐH��9L/GZ���A����f�Rb�'$f&�e��;2�Z��Ċ@j�o��䤣`]llQVSG���]��kL�e�4�,K�8/Y`Z�љ"��$��du����6�E��X�^�߅���S*'bD�ĳ*L��"Į�� QJ��ă�mC��,Q3�L����-��K5�[N�Y�������;%r�B��u���!�U<r�4����[VQ��3�V*zBe׻N2�)�$�>ou[c���x�N�<2b0\aj���+V�=�X&ލ���^"�� A�.@��y��e�߹@�5�LQt-{ ;~�Z;c\ �,�T�k"D���x�=�p�ub�Y\�[����;`�K���P�a1�E=HH�\8����IJ���>�8��ۮ���-jInW`rE�i2m�R�Г��+@$�#!#Zfx�U5U풘��%'v�_zs�C�2��˖n���e��*2������Zl�׮��䙓佒�x�=�#��nҺWZ �"��8i��&y��4#�A�B�{)��G�����Z�r�����"BL�.2�edH��-~���p�{�E�QXPe��3�I���l2��}��D������dN�����\D�@�G�14���x��_�?DA����ơ����o���!��2�]�xh��!�u�P7T�VB%���mkb�􊌀$���O��&�����ݤmR��n�?��c����b$�5u=��잭s����VXy�&�!�oj&U�d2��WX��j�n�ĖC6}�쮻h���-���MÍk�_�N�M��m�{n��=�õ'��FH�a�ø*@h[�{�l�la}do2F�9��=���Xkѧ��ɍ�"*2a�Z"B$�K���;�����&� mK�#.�q��Y�h�g�4�l=�=Y��wʘ���1g�"j�)hG��w��cL����Ƴu�<�x�#E-}_tk�"��j�s7M��y��2�^��dW��o�0�]��T�X��ۨ��#u �A��B��F�@�Ԑ4-50�4M6�*�UY�;.̶z��{3�8Q���;b�o}�[H)q���E�W��m[�����$�m��ZZ�`R�XO��%�Ih�h��c�m+��_�~g?����փ�4��5K�0ą�T��^(+��ޓ��s@�ʛ���T�\�Q���#xEYL����n��o���=�}��<��T�����k-'ݽ���p���$��Lrs2���5�H���GDG��o[޾��&��7Lt�)O6��4(�*cryTʌ"�>�����i.y��ܳ��T�P� Sj�y�AJ��K�}az1��#��m�#����^o�l!��y#�j|<���]F��ֲ��M)E��'������	d�\����=Mg�����z�WDL!(��(E�伏��x&<��u���l;������S�I1�$� ��q<�,y�v��cp4��w�|�UbϞ������_/�X-������Y᭥>w���8AR`�Pz7̼nB��CJ)�"I�c$>�.�Mn5���>�v�"e&*J����3�A��R���eڬ8�jT�#�	�u�A���NPj�q�s{ͤ$(���f��x~LY���WC�;�AU*�n��%E��Lf���b���b �u�k~��G|����д-Zk��9릥��ԓ9��!�C�<R�v"x�`{R�T�@�4Qp�������O&7�R��"�=/~�|�7��y���i��B���b2E���|�E�\D �v����ڎ��5]r��E�U8�6�~v�>d��'��b+2�!c���������� BOFl����!dA2,Hʀ)��b0B�u=��-]��mÝ�O��D��%M�R�j��PMJ�ȃ����C���?��?rB�#�B�O%B+�o;ʲĔS�����3wa 3�NL*���؄���11�k���}���V��������-��Kd� ��*��~(W����p�(rm��Q�E]!e�B�m��+�������?�o���]�(�����S��ѵH!�E��bR�C�C�F/��v��m>�����c�we��=I䚹�b �%��D;�8�K��1⑨� �h:O�9��`?n&1��������;2�`�¨��?��K>џ2?=�9iY-W���:I:%��4����\���P���ͳ磜�m;��%��3Y�Z^��pŎ{�C��mr+�H�F E��	.��sL�"�="�qx��j�E���2  �~� r�T���`߂��>�n;����xcBD�k;\�<�F!�:p����R�z�C�6�t��F�� 2g��Y��T��,$z(�D>�i �L𝨀P�����FbR(=d��{�В�;�?��۴��4pv����~<����[.���1�"�㤞qyyM�zN8:c{u��=�1�<d5�p̑��de�Bb�'OD��(���R	n��ygwd��:��n8�[7��RRY
SD�x'�li�EIYh
��RVS���j�ѓ�����Ft�a�\�����_���Ĵ�QV��5��i�p�3S�R�VP4�gZ��F���"N��K��g���,f����<9%\����1.��p�� ����%�m!Y&e�ݻwY[A�N6>1��#s[j��D������@��3�{�u��!г2
&���Ͽ��?�{uɳ����'.�u�NG�,LI��\���� R"�]��IY���?���0/KB��ڨp��Q^dq��O���x��9�7��
1�9�&��0)&xj�H����5��xg��Q��0Qc3�W(�6�xK�+DY��=�h��z5Ԕ#� �y2ü�|�)(��!13YDj���U"T&��H]��%݋�2�>��9�� �2P��%	�ZI����6h���w��ʜo[j$�2���]ܣ�P�(�)"<�g3�l�5��.x��m,��v�L���޷�	�ƄU޴5�-g�K�.s9d�!#_g���B��]�i-ރR��"�v;�����~��#�:�<)%b�5�B� ����~�[��{�}|���\���!�EA�ە!|�=B䎯$`bJ�۞��������uw�ك�h/�i�)�����p�l�� �x+��2��u>b�E��Ȁ�d�Y����vZ
rB�1��$�uwn��������)=�`%�jo�'�8�� ���ɳ�3+O+�	��e�A�hč��!E��N����B�Ā�B
*-(�>z$���^L�2>%U�CR�@\Dk�˚���KƎA��x�9<�} ���m���፨	hVW[�O<y|����,���v-Z�,��k$EFIf���}
��-�A�i ø[������+h�����cWk��ei���LgS֭�b����5�TS66�d����_�7L��	�:���_?cu~�zy�.�a��L�)Gu�駟�v+Jey��_�=�w[D�smE,	A�Y��ň(Kdi(JI*�\y�����������Q�����o��}O��.I��lY^��}�$��-o_C�k��t��	�� �#f��$�c}@y�	��S)MkĪ"M�S}|�O?�g<��3��Z���Q�3)��5������ӿ���xd�Ւ����NtM����G�ٟdb��+C�umR�$Qi.�)���㏙����	�,(s���<Yoy��K~��_���?P$��2e���bJ��Bi4.9"�թ@�4�R�q:��F�ɂ.r��.�ޱ��
��+Tt�Q�����prv�R��mpݖ3aI����c�4�8�R&KpAG���DV9�]����=FNJ�P�͆�v��15�j6�L�5k�x�	�$q�qG+U��B��P`�g}~ΉOL��h.�;G�J��q!Qb?�:���^{)�s۔ܮy��s��0H~K0J����[�F�VL?N��VHD2�����N����Z�p47��a�wm��E�����O�ō��Ӳb�o9}δ,xp�/S����o-�V$��l�Ȅ�3�03f���Ds��m-W-��rt�1��+l�����c�-������!
�Ȋx"�k�I�hߝ|����:�$��
��'��$+���J�����B7�7!!�6�۵����o��n��[���>I��z��1�6�$G.�T%U��*��#:zW�7�<,'&1�':��N}TlK�A߶�QdC9Fڷ��ߌ����я����k�sR�R�5���+s͝�ǘzB<*��@ȁd�"_HZ)�bp�v$U���j�Ӹ�c�o,������.�"3��I�m�)!���$m��c:��-ت�u�S���3�{�I�1��L�������I����⚫�u]3��f�t~�aK�Ͼy����)�d-)ee+L	1K&{�5�	w?�������S�L`��.Y2d������k�WW�޼��Oؾ���Ւ���A���J�,�+�3��I	�������>�������/�e��uH��I�����~��3���gǄg�������?���9��|��7Do3���\V��($R�и$R��=�ɟ�����<�-d
�!"�a�:�r��9��S~����o�}�o~��/-���'������6����6��)B��;��C�\1���ÿ��������%��
I��\.W�It�Rj�q!����Wt��m��d�O����Q%i?齣�Q��#�����?��_S(��;.߼�ճ߲�8'�	�Ԋ�rE���u���#�	��o���?c}�5V�sn�i�    IDATW�V	�Ȭ�<�r��SSNj�'��������R�1�n;�� 5�I�6�+9�v)���6xj�	� �DJ�"�<u�z:�m2BN2 ��>�1�Cۖ������>��e���(��K�B��t�m^?{�}��-���i��<�mW�չ�9�:yN�<ǋ��t\-��Ri�m�W_����=�<:)��#EJۻ�Ih�(��|B.���zt΁=���ho��B�{��.�\~�9=�n:z1�^���r�F��=�2�#��o���z������|�R��h��D�!���1	���Rj&�:�JچJdd
y�"��R�C��@o.�!���!�i	3��Rb��E�f��ٓ>C����G=�o�>D�	GZk�͖B̧s�W+�n���c�N�h޾�5��<%$q�#	����4 >��!d�E&&���鮞����f�����1N9"@HI��������u���=�Ŕy/���7/^���[�<¥@�%���v"��#�$Y�V\l�1*���rr$���L�*&%���Y*��y
�"i*US��mHF�./�lVL���@���2yK����k�tm��j�b�o���n���s��-G�r,{j�&H�TEn+R�")E���;Rs�<���.)gdY��Z&�A��h;ʺ 	����b��)�T��d�gϸ{�1o����%U5��m.��GZ�����t8�.hI%��ǜ޹��߷�JR	.P(K��;��b��>�����cI�{��o�ί��!(�'��c����h-U�)鈺§����Ϲ��?&	��j�7��~sN�mI�񑋠5]ױ�n�wv�lZr}�����"7�ʣ#����Y
[:!&�(�}bnf袠I��������	��q��g|��n��Y-�}�,'��-�d���9�(U��� �9�߾"YC(��e�]?:����V4L'�-z2ɶj�x��e������v��v8h+���;(I
-�r�u�3'H�s��6_"뼇�h��0�n@<3�J�Q��:�=����}�u�m�~��~P���-ᜄHb����Q���g���=}�G���xC8?�NQ�]2�bD�0&ϊ���3�r�Ń�z�˷�|��J�WK�H�mo�2YL!��
�@���m�(�F℈0ia���AnB��!~�w���)4�t. �Άy ��b>z�ȣc��RB���r��#l�C�|�Yj՘<&�0$$�!j���Y�D*f��K?d��Y�HSȈ��g֨��\��R!�����i4���;�.������������
!ax�p����v����DDD�0<v�"d�Zr�u�u8I���Z���)�4�E]�j���C�W�P!�E���c{E$�<)��
U�lm�������͜��!���)��KA�����O�P�ѶR�� %)cO2��&&.�Yƣ#ZUp��.R�Zx~�w�=�p��w�J�Z�(U喲�����;��]�����|���W�sG/f���,i����
��h7���P'������-��0I�r�%3~��o��'� R`ZN�6�At�z:��;D�'G\�K�4�=:��
��*���҅?���"-�P���.��� ����0;�<Y���5ǖZ$*�UDJY"D�N%R��\���7oIuIk�*h;�QU�Bз=����(g�'IU����g��,^��;�=��]����h%1�����5�+̤�~�=���5���Har���d=��LkC�m�T)�-�y�W���r2�	�������<���Cd�X�[֛+�m��-u9g�z�3l\D��ݒ�C	M;�!����P8b�;Q�d�uH똜�����_����bc-������k��h�}��v\�~���۞��^��,sڵ�6P���+Y҆��<*�(�H�5�����(�cJ����M���B�Y3���P!�A9-���c��%R���{OiJ&Rh(fU�O� M��%:����`��@bk;BLHS��m����;� Hd&�Ò�� ���ۊî�[�1��r�H��b�<@�S#��)��� 	�BԱ���%6<��g	��c)j��h�d−ii�����{<��t���BOX}sͯב�O�����~�5εԅ��,E�5R�	���*bt�%r� ""��C�p��rI0�('�#���@�@�d�ܫ�[�{�u�D��,��	�D��{�(v'���� �����Å3��k�c�`�`�C�	-c��W����c���Ū(5f *�4(�%����c�J��c!mL��߹�>�Q�mH�3p�v�K;h~�s�C˯U�]	��S���ۿ�&ӌPθ_ZgM���k&A3���\_�[���MӰ��p|z��M�o�dh�LȘ1\���ǝ�ᚾ��{����ˢF)�����0�w�r^O 6;�Ч�����]�8{xð�jWw����F���)�������dB
۷���rw�*~���x��ZD��
�%E]�3
r[�6�4���c �<)���	��f1�q����.d����AcU�)ɟ�ٟ�(���9_��>��v㌳��>�a^�}Ӣ� �<cT����\��Z^t�3���`ѪF��)3�����XKY�D"j`��c$�h�uD�~?vy�Nc��!���("���g=t� %��/�~6���3�� ��	�d�l^��畆���㻎iY�6=W��SЛ���I*�:C�z�t�TQx��!�������rͯ��'���?�(
Br�!X��̄ �]*��+�?N�ZS*�����k�ٔm�!��c��Sp�8F�%FJ��Y��m�=\��{�Iɶ�6��B
��$��-ۻ�'rh�REFLb@h�TYs]*I5�P���M���a��.��C�(��w����0f��ux`�RN#7�����v;���%���!r͞�DD�">$6�o���'�������E�SA<Hh��"d�3��dTb�M���򊢔|��N�NY�}Eg{����p$���r�͵�;;:&Epӿ��R�A�蠇>�]�N�{6��>C��ln?v�����b��}� �����Ic1b�Ç�JٰB�ɇ<�@J&e�G؊uŰ?I
5��r�PX/i�〚xc�/����,��9�<q�9�P��Ϗ��}��p=�L��$��v�fuq�����	zRq�l1RO*|�fH��3tB�HYj#��zSZ�9���;�w���~�����V����ݽ�(��i�ێ�uĶ��^�˟�� �S� ��(�A堇�׬�T,3�u�&��w���R�Z����W�W��l�֚�O����Xm�\_]f�y���)D겢�sf=_�8;;&i��J�H�Ȋ"
��3��9hN8�}�s�-������(�����Wר���2�I8�p����G��⚖�i��C$�=��p����r�X99f:;E�	R(YF(rqq��_}��jw�B���m&�f��a��!+!�GL	;�s��Xkw�)e�l2�k[�..y��%Z*@дĈ6��(X�fܽs���ɰEQP�3�lʝO?��GO(�D5%ױ���kX]������.�$.߼�?�{��5��EQ�;Bh@�`z�����<�{�RI���~��fF���m	}���R(�s��͖�oRX��� ��9{t�{O!
MY�7�!�w�ڡ��wZ'R�)�싲.s@@n�;xS?��c�M�x���%��Vߴoc87�ﶝx�?��m}��9����#)���L)��f����._�eq���.��G��cIO`h?�߀R���Fbd@F������o�����:����c;��w�N��sr��U�����	��-�j��#�~Hp3�9�qg~�A��3�sVW�5�,�|��ټ�*׸� �(�Q3�M�� Dv�r62
)��7-�mO1|��>n��y���Lt13�%H%��[����=<?�[��=7.b!K������8����O鼧���S����(�k��ZG*(�@�1J��Z;G�k�L����~F��Q�z<���)Q*���ܪ�m�ۆ�.�\^�6�m*�>�EBi��F%��є���{���uȘXTN�����*0�c��`�-�8Y,8>>bq�������_ `82���$��8�|Vqz�����$�"��SL��sp�o����
)�ُ���ϙ���+��� 8�����"��S۶tmK��ҵ-��aF<�p+RQMg��"�2E�vKL��z���k���k�qͳ��RC�w����+���{ 	�$h=��3"�X��ƴ�-�e�ʟ��3TT�d�>���z��b�R���0����Gs�s6�����v���B���:E�m9)$G���0_Ly��	'�)��)�,J$2�C¹�S��u���5�v�!���|��WІ�oi6��͊�K����>�Z���-�6�"��:|Hh���O�>壏��R��R�RZ:\��#���?���x��Z0�M���8t$�DFBc@���D�,�((�
g�M���ɏ���(�ly�۶���;�W��c�I ���
z���` YJc�F%m�7��-�O�=z���}Z!�b�І�4��׹��t¨Di�("2yf�
��_���۷���=oD���������g���}(���}�q��E<��Cȡ�^AP w�����������v�u�:�R�$&�ط*�^�E'n���<�]fG���!
NBJ	$���s�}&�	%A���}�vJb��9e��C#}��t;H���m��>�^`p��}I1�nFk��4���/�`]�΃��bմ�� ���C�-���FE�Bb�0J%z�0Nq�.�Cp�Û~���2A"z�
BRO��E��n9�O3�9F�͚��,�m򻵑0@l�H�)'H�ض6�	�uD�2ۘ��tƴ��]����,�oQ�SO
�fó��z��C�v8�e��88w2O6L)���}��z�횮Yg(;�GJJ�	�.�VJ�v��j�������5�1\^^Y�'t�d����hZ�2���Np)OIL��K	)9Rr�ǔ��m�!K�]��cZOX^]Fgi�[���"��x�Ѭ7�	��#�1�R�i_�{5�3A�ZKi���jKsu�S�$E|��UI�ni7[�1���4R��9ǅB\���xM�a.I��N)95�ޒ����R+��6̎�|��G����������uv�)	�B猽w4M��޻���%�z�k;���eH y��;���z�p�� ʒb1er4G�{���=���@�˟��_��g�R3�j8�2�ޑ���f̳D�*e�KN���V���EJ�8�$H�ǯ�=]�H1��ލ�=�u~8X�]{v[|�]�������r��|�f�F���(��I�䫟��|���''\�����w})�@> Sv����'%r�5�Ɍ��s�m�S�o���)�'�{(�@s��o�>��p��08w�h��_i���w��bh��g��?�[N�m���ُ�ޜs�.��$���d&20�!��&�t#J!�0�G���{z�lDHM������È��!@>Y�'?�'�	���#���A{�a���;n��m���};�g(�`�S���uù<|x�ӳ���,�*]  c�R�]Ғ����z�bȣvo�/��:��fT���ٱg1��HC��)�B#b�Ԇ�ݢN�a8����RF	i/�f�
�u=�u��6Ȯ%G!:	RH4��zu�st|�Z����1���C�e��a�zK�;�l�tyr�NU��#�����"!$�ϝ�}ߣG�r�G�"&R���Qx
)�#c�.�fn�T���x�cV��$Z]������
�3�r�����$p�%Ȕ���%u�VtJ�vH���<�Q!�F�T�}��;��΅!,N�8��3	w�n-�Z!�P+RVg��c�f1����k>:;&�G���v�v�$�!$>�sYMi6+қs�;O��,j����_p��0�'\.��|Kg��ח�c}}��/_pr�>E5=hN� ��r�2xCr���5���m)w|&��.+��	��w�>�4��YD($
c�R�Nۡ���D�"�1R�-oe���-� zXʺ�,2�d�>￼�5"g]�к�����x�KB�]S�m�	�t���}���]�ۈْ�6�}��}�q�EH1LY=��?J)�fë/���b��!�h֯�0�rR��#�U�ȃv�Q�!�h$5�S|ʭ��CƄ@#�H���m$�}�)��Y梉�Ba�W��ރ�|���������j4.��pH����݄'���� ��l$ E�ഄX�(L��a4�z�m���d�� �3@�Ch飠�z�A�n�o�!�X��&�.�MG-���nrv�,�%�ݮ�v�����(j�q�og�q?�QJI�j�����7<|r���)W�m��3Lk�$�����4O�o	z)�d��C��|��}Mc������X�0�%��1RC�Uɫ՚��C|�Tu��(�R�g�H��O��έD�bq��蘵�XR��ozʔP�������7��:�M8ټ~�-�`��u
�53��ڎD���Kp�~pmC�Y��훖�uTJ�i�6%�,�����R ���k-�Z��hY�]o0m�qa�R�wB+
m�6����'�h]Ć�]P��ೞ�(#P6�ҡNC6�j ��h����-��cJcr��qXQq��R�D���[���Fda�}x">8���ux��*�i�{.�r����z=vr��A	޼}����(�"ؑ�Yo&e�f�aڵL$��������ÿ�P�
�}�wR� �������%b�i���Čݦ)�'��"�]�ؘ!R#�'j�p*C��PH	ۦ�K��q��ﱸ{ƫ翡�l��#�B�S@��Y�mD����x��F��,%Z*J���]�)L5���՘�t��|Ht���I(�t#b�^�{?�(9��(��>�
�w
�A҇l���!2��[���`@�w�����$o9==e�v���s>��NO�rѶX�bb��>)č3��ZKdXk�&�����k��f�י+!n��b��DN^��8���[���Iʛ������UɧC}�y\����܂Q���j*;�!��J_<�	;�=Ȯ-��2��ߵp�7~O���N�Ć��i炜�Q2R�����Ma�ß��;!ҍ�rB������y;|����]��̢ۤF���%���2j����Ͷ���,N��y�v�$���9XP�H��(%F�!ɜ���~��ǃ��qw���򽏂2&C\b��zuj!�h�t�ủl��O���]g�Vr��4�d7IPO�ܹ\�E״l6�x@-��hN�M� �!�	-IIl̰������ч<��(ݖh=M�ж-�v���[��)��~{N}E�=��%�u��!R@Ę���׳4����ftmK�u�bʝ;g��(�!�Y����E����v�D]TP��.d��ii�H��Cq*䠅�;Tz�ج�\_^q�{�)��8��5)�����n��(P��}�z�u���-%�l ḘT��BӇt�<2��ȃ�r��ry���c^>�����	�,��P̎�	�5��)�A���_=�ُ~N�$Rz>��ӂ���YR�
����L&8kѦ�����L|LtQ����c�D�%U��	M38�@�w�q����;�횯^���L�Ɛ���jP�|檤@+"Y�@Hq�Jc��H��dF�
�k��SփWJ��'C�R��тmے�Қ0�T�QN{g�>�����[�A`�H����~�v�I��{�{�������-����>���ݻ���|���hJ�Ӕ�K��h�����p����Y�>΁��e����}�o�2ȉV��Y�)"Y�̆t���W�A=mX2u��_��2�{.fr]�h���)	�'&�4Y�6Az���uL��f����l۞���"�J%x�}"&� R&�)��O���T�Q�Y�B�ʭ1>�u]�p�Ph�3���;��c�2F���/���o�[n;dT�"��$%	:k�'5��8|>N)�nz�+�����W�h��V|IV���$��L��b    IDATd�Թ��ؑy$*kR�Z�BH���Ie�b@�P��`S@�@�JKZ+�������۷T�N�@�X����놯���/������1���O>�;g,�|FstD��K��>���������S����5�m����+��t��\��K��j��	W>Ҭ�h�@���d�ݳ;|���|��g<z����Z��!�>&T6�5��mRe����&tE�.A:���v$�fbWy����mt��3LQ@'���m0fʀ(�f'�r��1jv����)�r=O��m�O�.Ydt-�È<+��=1X���Ϟ��^RΠm8�tĤp.z
��E������"
Xy�� qi�"���$")�r��z֛+"���r�+f��׫f>ϓ��۞�r�O~�3^�|MksO����(4!v�&R�D������"��2�v+b!H:"cC��.0iʝ�ߥ�
S������c�\.�h��T��Bj������$%22��Qx/�'���L���+��U�O��dZ����E�*80뭵�2��A���0*�%��p��!����aQ+�"Z-J@�&J�����@W5C�����́�I	3��;�02ە �L\�;�8���0s�#�)# ��C�����1d�	�y�1����@�m���LHR���"�����_�|uű��ꊠ%^F�� �\0�4�*5A�u ?@��ID\ $*E)�ޤ�L������G������8?�y�p
�|F�\��yA"�BN^����v I�ah[��[��ZLh�P�!�����y�XPv����f��sۡ���v�|�)�vБY���co;Xd�v�B&�;&�'���r-s_O�ؾFr�χY���o������o�7C�z�n�6��3?cv�p�4�~����svvF����-����2�)]�>O�����#����51L�I"S��H��� �A��λ�Ze6��[\ہI&�@�����)(�F ��K����jŋ/x�����jE�4���<��������/'S�Ն�:t�v�Rc���;.^�]�*']�J�����js�1��1�`(Y�1z��X�6l��T��9��?�C�N�s��_�r�K��9gc��ƛ�9����.�	�{�j]�|Oe� ��a�ZE�dRq||��-9��x{��K��Y�N�y1�l,��I	eJ֭E��==A�Vr�@�pY'��ϑc�a.uY��� �9�L��a�7xGg[B�TU�y���ꊙ8���w?壏���4?�я��|���Ȥ��ȨKӵY	OJ&��������1�������Z c�]OF�����c���k�$�)sBr\�=�_|A��;������;��]ǫ����g�MGH���"��(*�
��j�WW+�|������?��w��	�7k�ߒDĤ�kW�mƿC uVv��"�;Li�͐���>"�CYgxc����:1ח��g��-Ю����{M���{/|��8@�����6�}����BbL�$�s}yI�\3�̐^�w�v�u��:���Jc9f,�J!d\f�ܔ�AI�ᑥ��;�����xB��sT̏�\]]��@uim�?uxl�3��{|2WI���q�!E��v�=$|���bpD�P���+��H9
�ffo%�n���͟�IA��v�ޮ;�7�~����C��s���q���6���w*QJ�u��CEx��.���/i��P��r�H	)�!_6"	4Q�(��bh9i`�Ɣ���s�ܷ�ŘKB��Q>d�Zo���%G�W�<G߉L�36H���?h����d��	k-���3����w���~�O~�K�vÝɜ���ѭ�\O���Q�����b~J*g,��GǜM�D)��������eCIdzV�5���˫s���q��$-�Js��#�?z���=8���Gތ�q�rpҩ	!s�4U��j�,�9[�)�!�!ͤ����iX��xow(�f{��z��*��3_|��i$�n�d��]�%�����7�%����=�p�̼y�*VY�H��D�(���ڍF����@��0�����n�b��*S�HYŢ�Xwʛ�7�Þ�aGĉs�䭲�(d��8q"v�ر�w��.�lږm[���	Yn�l�l*�XhĚ���uӰ\.Y.��3����������M��>����K�7���"�-:�~�hf�)m4�M���|u�������y%�����яy��E�=����Y>!Ӛ�(���!��&F��seB�t�;���p>�r�Do^p����>C��l�8�l욯����4�%.颤n>��'|��߲���ưX���+?|ȣ'_AZ���?'f%�E���n[�4d�%�u��l�l+��?��ι9D�c��Q��������i3u�LD8��]h�i��6��%��r`�qt�9�p>��6�H�d�]�K�
�s6R[s�5xD"�ܛ��1#�pߡ�;��?�R�R"�!��M�02!���%��XF��{���U7��q�HD@ң=��][���5���Ĺ�Yua/�{���a(1��؏9��� n/�n`_Y���iP�����[�v��MR�w�1��:C��J�kv�xB�A#���u̲;����7��@�c�U]�tx�c�h��{uq�҂�LY��:�)+Z��t���QRPf��$ p"y�1*�JFH�:�G(d
�R�s)��=� S��Pp:�"�K�2�Ŷe�6��Qw��E�3�LY��ԛ-JJl�R������eL�k�^	2fbmj�iC�"�Yɬ��N朝ާ8�ǫf����C^��/�y�⤜�����8�q>rqu�v�AH�7dA��Y&~��R)�^'�օDIk�F�Ny�-�����d�)+븾x�˧����K���"��j�a�޲��4Mӭ˴~����i�O��ڣG�gPe��3lt�F�w�C)�?&fD]�(�Ѻ�|����_c�4/��H]5�#�n����YK���r�w��u��W5,�.AF���.���:�4�m[jo�F��O�~��|�BAuˏ�c>��246l�e��Po�e�1r2/89��MB�a���ж�f���$ţ�L�z���P��IA�|RT`~:#���7/>�?��G|�˿E���MU%���C�S̓I�÷�e��S��-1(���j*�&CǄl�|�Ͽ�/y���bM19�!��Y�O�O^��:i�#S�TtL�%�I����چ<��Y�P��xJ�;��%����L��(6���c%�����m_$��s��/:�s�������J�J�F�P,)��L�c�~8o��eg�����B@��ف[j�����4*Igv�K�����[|E"9��Q*�~� ��AG1��w�Tr�6V�T�b<NĀ�@�׻.�(j��~o �Y�PQ�qW*1�a�{�u�D�cA�`e&D�3�1���s�l�Z�Ǭ���~;�&��E��;|6:vl�Ǯ�ZJI�5�0�W�.i\Óws����k|S3��8R\W2H�J��B+S�#��0��4v�#�5F���̤�p�Sh�4dENP��#���M�rM;=Ad9���QUV�,�R�v�f��2�L �[Ke-�����s����F�5�����nȳD^p�Z�}��	O�ݰ��|�=|1��T,�	Z�F�#A���3���� �ٌ��׼ڪ�WU�pP/#J
\W����BL�p�łZ>C=z{�O�է|~u�G��v�_"��'T�G(Mk=U�e�F:�α�EvkAt�ф���l�H2�j�j�B�	�(E��6)g�:|�ȏ����e��X�ߠmCX����iۚ�l�2k�@�-ѧ���fC4LJ|S���?��1�����>��r:ek#H�rP�Mے�"q��T�S����OɊ���l�'3
#^��ɦ%�ed�)�r����O�����5�bC���:�/j���L5M��5�f������cb�T�E)E�e0��4���3>��c�k�;��NOR�h�Q1�[O�%C(ʣސ���(
�ɼ$S��i	�v���`�%�{�S������ܫK8N�(�Z쮻�Ab�ý�ۏ�.��'�������
��{J>&�C�>�;���{�kғ��0�w�c8�o���	1t�=*�}:=��%Do����>�O��{H�	�H��v9�!бi)��cu�BO��{����F��$����n� {Xe���ev�L���ޫ"q��7��g�o��Z�����[�����`J��l�c�x<'�^�]�cǏ��.xjoW���{C����C�^@�39�+�
��b�Қ��~Ľ�OX�\��n0"�|
)�rW%��|�:�%1&�8�y���yچ�����=�s)�Nk��("�k��-��Z��5��9.WXkɵ�78�w��r�����)%��H��Y�-����v�^5LN��Īa4��)�G|/onX7-�����@�x���wp��U�^��U3��&�3�優C���	Ֆ�nh*��`\D6n�b(Bg$��h���!7�����i����Yf���Ƿ^.��x#�(��N��t�]pm�5h=Å�ń�|`�15ֈ�$izrB~rB�ג��z�6-�zդ7O�4��s�;'{���ϯ�.`72�1>����R*�&t�LD&ڠ���%5�I���5W}���klUS�L�����r���L���M��(6J�ԕdBP���f�馢i,S�y��]%�2)���4��������g/Y_���j�ܔ�(�23��Mǅ !��A)���9EYRw�􄴾��lZR�KL�@F\���L�6V�G�����&�u�n�d��ͤ�ZG�KN�r#��ں!Ӻ[rp�B";��m]R�A!7I��{��NEBVw�hO��!�Zq�����y� ���\���vw �	%��U`o���C^��i�wv��B�;�(�HY�C�C��QY�L%�Cǿ�P�����������<��,��a�+�8�קb���Gb9��.��{�R)5B���/&Cv$."y)c�A��튘2���O(�:��W^��F5�����w􊵟�c����w-����F�x~w�V�q���\;O~<����y����� y�+�(�g�l�9zf]-��.�A.}�i��tp]jH�A���|�"%���Q��G8𭥩S��sZ��'%���o�Je�zq�</��Yܿ��<m�%��4���������k��Эg&����]y��g�^���ez�Zb�'7=U�ٜ�,ȍF+sBY�I��<`:����l6�t~�f񚥵�\]�o��*5�S@�@�)J�#6W��U���=�����*Qk�˖i9#@ph��g�</��Ȳ��҉E)�m����U�g"d�1x��H�	����1���? /Jd���:	
��&4�x���կǉ*~I}�%�5��SNfsژ*1�Q��mKS���FI��z�u`]"�i[V��o��缼��ZI�sN�N���m�P�53����Ֆ��k^^\�`������(���U��WW4�W���ۆ�e�|�=���X�%mk��kT��1�%�����	m
�����Tb�J�CCnJd&���FK�f�rI+*L(Uö^`Q�T��8v��2�;2)rC���m�mcǵ�1�I�<�æ�<~���ߞ�vLN��*���|;��}�����><(��w��kd8t(�(y\tl|J��١�1�xS�Y�1&߳�a����p��N/���	��.DJpD�K�;fpDF��봚�3��fE6)�*����\�܆���C�N���R����z�cKR��ir�	��!����q�xb��?�h�FHM���>��{����1����˫�� i�АhI��s(�1i����������[�<��[oᯮ:�� 1t/�B��@H��V#Rݽ�R�ҋ!|����E� $:&>o�RM�V�LiTH�MUD��������l��ų?��-QFj`�^#�����E1�L��r��}�1�j�Dg7�T����Bi]�g��B�.
|k�e�TGTtDA0�
L�Y�T;�X�m=�>�y�ki���4e�%��ۊ�jö��&%a��9G�G�.I�dYk�ֱ٬�������|�O�~Φ��'o!LN���1���sTR UA����(d`�Z�Y��G�9Zv`�lB��w�E�.QgB��M����V]�d�(-�:�s)iS%H]60�	����VK��Q)�tFM��m�i��Ȕ��-�՚ɓGܸ��d���qZk�<y���^E��ε�7�_/��H]�x���1&!�1�M���򊋋�"*I����Q��>2�L��-2j�������\G�ct�1������S
�:�a�֊,��%_f���*�<��X	N<*7�m��dG��ؿC�ՔeA�i\��چ<�PBSW�F���+���^>4MK��JZ��ܧ���Bo�����>�ǹR���ɺ#���q۸9�}J:la��1�z���S���I��� ,�D����=������Q��z��x��ј��m1 �R�􌀾L1�H�a��&v�9��ίk�2�9mW�!y�=�o�!��M�[���<8ߒE*Q���I�D�ZQQ%O=8�R(����J�@"���Q��%iZG�$6ơ�R��!;�g����F��H��O;F��=L�~�S��cJ��&����LG�c�t��6�4~0Z�@;�;�]1��8��x�&Ϻ֍m�6)�\-y^{�߿��M�.W�()�I�Tf�K�LsJE��
Ik1�7M�]��)F "P��9����|����:���'|�'BY��cW�T���%��Ͳ8�,7X���lZ�y��(Dǉ0�8  ՜"Zdgӌ��E���Xoh�S�ʱ!��^N�ْjY#���P8�Pq���-�O�4V�8IU׈��qR*�c$TJ�+M6��P��'�-m�����p��cB�i�B���ׯp�3�́U�Ӓ���;���w�Fݬ�<�`�$QE�:y�!zZ���DC���"'/��9r�b�n&�f���	���ٮ���2��l,˟o5���
VFb��8%�G�;C�%)�kJ��Nz�R�-Mf�Q���ak�2�Ef"k�F�H^��l�(�tL�@�$O���lj�?9��3�UŢ]Rdڶe��R�5ֶ�M�vQq-+��kB�D�|RrY5�	:x����S)9���e� ��8�b��G�N����tJ�gSW�uŢu(-�����m����u[D�`"TkNf3|nX�����4d�!�9	ѬYǈbFnQ'�,ˈ1�Chߵ��T��'���t�o#.ڄ��5�
�B(�����
�"�D��V�J�H��X^2�)(y@{UvIbc�­�d`/�����ϳ��O�}�<��$"xB�!-$GE��,�Z��mED��M��#�j��z�h)"���"�Ó(	
�� �2�:J$���ɘh�{#�CJeb��c����Sސ�g4ZQ�����M�-��{��&'����}�����҅�m�?���[������{�`�C�c+�.x�������	���K�Lc���q|_��m;<���4���<x뜓��^�����
���u��N��+ A�h��2�&v���5��DE�]����_��3��_��=>��������7-�"��Oy��!�W�M���R×���DB"�>ŝ��N}�Uj43՚�sl?�����=�����O���{��l=�?�3��W<��ԫ%:7��z˛�HBa��R�̠����3Ĺ�A(���i1��dN���g|�o��-"��ϯy��{\-.�ş�9~��D�hچ�R����ſe�z�,+P&�:v(W��UGb��'E�
-�Θ���g|����=��q��	r[���3�j�p�ZO�����2	Ā&t9.N�"u�Ӑ��|�Z����B���Z�<��b:czZ"g%Z*~��&f��wߢ~����0:ps}��������
�'���D(SUuSB�(M�Fih�4y"7��d��'<</yx��i0��������Z��I�T���
U�M�:Z��Bmq�u��>e�^�� ��    IDATDT�,�k�2gu�����������/��k�T(bg$��c�*�R�,7Hqm���I�Sd�#p�v�3}��(bbI<!!�d��ZfO���{�ۗ�Qǎ�q��0�a�)�����9�������[���/��@*M�������R�H���^�������D�c��c�~��=s!����]춢�K��'n�7��F���bA�R00���sS����;hl<���z�:X7"Iq��E��z�֏�и8���ݺ�����H��S�{�J����)�`�ZB���a�p�ի��ӕ,jV��A�d@w%�.@����.vI!RDN����������Gq�ל�����e
2�������%���9W�6qo���<DW���Os��h	y�'p��r�ӟ�/�'���xu}���}N�S^=��|��O�"c��heM�h�0�(0Ju4�b(���χ0F`ʌ̗�k��-&������o��!���/��}�f}Ë�~�Z�FwIQy��u�O������ɻ_�[����EA���.�Z��us!��,EG�.QLu�������ɇ�P].y��-|ky���kf�$�Q{ANK��&;@�=ƀ$
BD_]�t(�J��8��i#�����'����?'�{��Bj�^]�\/U��rA��Y/	ŌLJ�I��V\��`[D�>Z�����9T���&È�}����	�~���92;��-��
�|�q��H}�Cŀ��"��RۆƷ� 9�\jT��C��90��,JJXHI&=/>���O�����FI>��_��?�K��F>4�RDRV����'�&*A���hA^�`���}흢�}rL�"���B���(�S�����;�&����"�
�샇}��v\��w�y��;��2�M�u��T�����Xq�QỶ\��>v1IY�����v�(JЕ,���T����ޅ�8C<�u⸖�e����m���]��a_���}l�!.�Q(��N�1��.��y�d�.�c����_����:'��|�6���x-!8�b�l���y��U�ｧ^�\\\3?���'�;�-�K���]�A��-�4�؂�b"FY� �킓�s�vI�Zs�2#�G�M��kɐ�ơCoz�b��f��[�J+E���-궩��V��B3/&�H�����͊)
�]��jCY�<*�Ę�@8Op�=�K4k�L�:~���nw�gd�Y�.3�JU��9�����������zAn�Kd�&S�*�*gY�=�uLL�,2P�YJ�� �LLto��Вe�#*�t:e"����◄mâ�Q�5�U<:�a�b�mqD�X,���Ti�ϭIJp�F=1&/�8R���B1��抧?�2D�I�N$_��o��xu�@�����,n��>)ܼ�1�h-�uC%*tH����G�1$jT)&sb`X��ŏ?��O�!3��3��nyCV��jE"��#0R��NpkL9VJ�(����	��OJ�Q��&55ɔ$����?Z<�g%���`a����Pyt�6�x�֑i�tR��@��#����
%p�ln�DŶq4�A�&(��(S�����j����׍'v���8 vyE�Cv�"����ߴ,�o�
B܃�s�?T�DG,���;����5���u���5��>R���^�*���!g�0H���s�zJ�~��6��؃��з��8$��C��������1��K�8������A0�Q��$��`��������5�nV��.���>���?��/��!1q��=8ϗ�<�4�/
-�����u��R�����%۪��WQ�9��X�(���#=G�e�֗ 
I���� x:�� $��加5�yI�u]�Ʒ�Z����9�2h���Zk�XL�S���]����a�Kr����d�:l��eDx�4�6LT�6��R2)��&yJB��3�y+�����������ʇ�9ND�"7��iIlk�匛����"�WWiz��l��S��V)l)�'ejHԽ���wDJ,�]s"RK������m��e�tY����[��1Y�r5��H��yB��"�sR0ƈ4��REDh����im�(x�4Lb�m�4�M���2���@w<ݵk�N@��,A������JƦ ����`c@��4���lj�ߢ��][r�RQ�(�;D�萤�Z*�L�7�4�c�ޑpU�q��n�%�lB���P�z�j�����sN�f�=�[+
	]3E����~e�d��L�#d2,;�)�cF�7#"5^r�<�F�]?yѵ������[rr�C����)��N����;�.�����і�c=��]��y�n=*O��������>�.�g9t;�b����}�0�c{�a����3&z�Ůڭ�njw�nV�T���G�758�PP ��uTw?�<�;���|��������qb�Vt4�2e�
��R�� ��ԝ���u���/�I�=Xo��Kw����>c3�⾵�������>�n�Yj���X!GQ8�X\/89�`�)�S|�����=*��Gr) �K/CD�c"Px�⤱+��.���"'&5Ԑѧ��R&ӂf��[{Z�ߛw$B���Dl4�ac@�"���Ȑ(����?D��c��v�����:5[���y�1�Zk�N�7����d$j��
雔!m�B�H�۪E	IUUH-Si��̦
���A�Ԓ��ydc�[�����ij���5X_SxK���� �L�c�jjB$�!ĈRI�)���d)�q�y��#��r�JcLa8�	�T��-�@��6�ˌ�/�B����\^�����\�T��ݟ�mAz�����F��O�^��8�P���y0(�w!k9�
d����Y�PGA��N�#���n���8�y6��ic�%�m<�j�L"��LsEK�]/Qn�=3�Y/�R:V_�k�r�|2%�"��������"�����_/MF��ԍ#�� �9b�8�&�9,�}rL.�)�o�ɏ�+�H%����~'٥��_E���A��돢��������y�S֏rt��{��њ�!�#����#����M �����(pJiD��.RJ�L�!�[��.��>��b�c���$����1{7"Q�+���,���<\��!=�n�{f��|�#F���/=N2^D�����uxܱ�1��У������5ֻ��eb���Q�;�1JѶ���KB<����I���LI�PB�@LW�S�9-Ơ4>?AvlyR!���+T�1F�4��\e����	��;��&��c����P�*	!��A!�EI�1�V�1d°�cr���%�v�Z��B�h��1�p�"�[����R�ZKvR&�}��s��l�׌wh!>:΀���d
a��5���iBde�}����zb)A�^lȤ��4��8��C���y��BK����V�J�V�u?��1��LkX�{���"E���=6's�%�����r6a�=��ݯ�������Tֳ�Td��	"�PY�}���+	S"��y*�:��9�4x'R#U -�O�*�QX�֨��4%�!>FHbDEʦ�J��Bh!НG�t��تAKM0>5=:+q�!m�a��b��	�2#����m�����ݻ:~������ZX��5��z;�j,;���v����ݱg +c�;h|��1ǹ��<�=G+��B<r�� 9v��(�NǇ[̥�y�b�Ӈ��Ů������L?v��k�Dj2�T�'b =�6�?�	y�|Kq�Ѥ����{�J;�7�Ĩ�aS�z��8;6 ��=E�{##����{�ͭ�s�~�c{hl��I9_��-���ޤ˿�Acb��'������7TUŴ�Q�)������9����c*�]xG���C��I��}�OL�T�I�l2O�W���٤d��DK
/e���jj|�)�!�@�c��tvs��оAi�$�X1!` ����2x�wg)sM^NX�6�̌`��q�4���1`�D@��H�1�=h���f�S�u�TL��LHp�IVR�nyB3�Ld�=���"������M��t!6Ij��T$ ��HyD�V�<BPSOsE@ɈV:�w��BI\��@�ƃ�2x�GF9$q�%~=���$���!b$�K��z�V�QeLb��)|b��^��+N�)�vd�lP��{P%^$tE�r':�R���#�@Y�iв@��!��"C�i�}E��9��\��PM�H�f��:�#Z�{�����׵��D���l�y��L��H$A�!:;���.%
���ӓ	1:���d��]����	�B`��RB�P':D�A����ҏ�ʨ�X��eS_��[<x�c��:��+�-+��|;���s9������Ȏ�-��~�{�J��8ܿs����1!����>�oD��zSj�"��*�$4�Ӈ�i=�I�*���w�i��PbG~3xx��(DJ���u� �d!E��|4�F��.PB�D���.��H4Z�ă:�A)3��إ@h��>�ej4	�uaR� 	�%��v�K�Cҝt�[~�p�1!A�,V+�P��Tr��� 0�.��p���{�iğ�%��Jއ�?rZ(I�wٺ]�|.'�<�\��,/��&r~~o=f���y
!���z:IM9����TĔi<��4>�x�2���lM]�0��vI���)|��+�lNn2��%��e[�n�A��.��?O��QG���f��^�����2z�*�1�6��ȶ�"2��5�e�L*�T:�2A"2��I�QvU]$D*'N%���H���<��L�M��y�^T�L5H�-���x6I���.9}����҈D�����(�ᢃ̠�[! �ilˤ�t�Ll��[b�h�m@��Vj�Q�˹�-y���W�%JC��X�z�TIF�Jn�g�)l[V7�xv��M� "k���� =eVR����/VL��v5�Ո�)y�DO�6�6�6��8Kf&@@��Z��&��!"|Hmg��SE���������O"S��CNr6���|�j<4.VĶA�	����k�&���w8!P��V��$�f3\m�L5NoQ����׋�m����7�bRҶ-�PXg)�%FT����iȤA뮕n "Bk�h�#*�V��F����]�M�|&*A�p��p�h\]6>;��vhꡂ~�HN[�9���H�aܡ
K���n�L��١���$���v���D��H;F�����D�ߡFr6t5�R*Z_���xD�h��z&�A
1��O���B9��� O��Tw)9)q��h�gB��`�۴��F�4	]"%&�ΰ2H��>�>w�D�1��ᡱo�ܵ ޴�ù#�,�@�2��踳Pb�����[>=
Ez�����-Ҋ�Ф=�B�p�������oh6q$���?�'}x���6x�_pLo��c��on8�͙��Q]��m���p������SDߋ@KEa��*��EE5�ȓ{�D�T�,BV���ٔ�������
��u�Wk���K�V�q��J"uɫ��DךVA�D�+��HM1�qM*y;�ϰۚ�h��\y�[ǩ�h#,������0'֦�����5�1�-����$\���Bf�Ep^��)�T��<+p�Ѵ�G�Q��b�$�-�k_g�6��LJE������f����u�@h9ӆ��m�Tf#&D�!���\E���2�������g֒�&�M�4
+,>��9��.Rd9��K�a�E�o�Qi#�mɄ&��&��D@ʖB(��)����.�dŔ��i�&q�M]o��Ln�FI�6������'�
E�����	�����B#
dVb��Tf
������F���|��-���q�M�p2+(���xV�b~:EIC��2U�:khs�|2Aw� *z�&��,���h�y�>�	��hˈ�I�)�Zムi,��%�¾=�y��ʠZG�6�⨛��p�l;4
��:���G����E���|������4��F٘��wc���#�>���Sw�C�?�]�+!}��!Rpk��Hzp0��@7�(S�T�	v��C����H�� uq[����I1(e{���E�{½U6<�>i�﹜�	�ւƋ�]��xBc�,ܚ���{��_��,��p�n���ۡ��w�g�Ѐ94T`Gpa�e�Z���޽S�	\_�d�l�j�4]ן��� S�q�=�7����÷��?D��X^\��O�����@��N5[�6�O�����V5:���(%�ۦi�1R5ujz�-���r��b �)��8y����D��a�4�OY}�&mLge)f3N��BrysC;�3=?���dʼ F���Uk��u�C5*֗��5�jhaXf9"��Ea&��Q�9�fCռ�8<s9�r]1y�-����kϺ���9h��g��ڵ�X�S�)�����5eY�I�k+�6A�.׬E��Z"��]�7�|���eK��ט��/�K�B�"%;�!b�*%oFOӤ2.D@��
�)"jj�d��͒lr�kk2��(��-�	|�Fi�uͣ�@���F�Uæ�	Z�],������%u�R��dдL�r�I�#V�l�g�6
�da%�s����D���q��Y�&U#�j���i�V+�\�L�H�����}��fL����z*0u`�x&�����cJ���V�%��e�!���)�Gt]�b�C�9��*f��4�������3�A���~�{�g��<�/��u��c���Կ��IQ����_Ӷ���$]ö�<�bJ��a�����F���0�w�X����w����x��񶗝1(�;�6	]�h��0�&1߉a��1$ �I	/����:�(��D�ؕ~����*�o�ЍW�M^С�vh�zӇ��g�hٷ^��w6Gr��s�uoo����B<�V�s�h^��狋������9y���������儺�'H��		Fu�]N������|�����X9~�k~���(�1�Q[������۬_/?�a2���o���Ǐ999I�V�\^^��石Z����z����)Mki�%�w��η��ߥ9?#WW���a���o�5W�����,6��	*�R�����o�=�҈n9�*�Gm���P�������ǟ�]Z^˗��	[+��������\����(g�ُ������(�[��t������]����?�����o_�b���Pf9�z�bq�B�ԉ�TY��s �M��놪����ۼ��;��̦%�5���'\��'��|dmk������x�ۿ�����WV�5RG��x��?��M���?�O�7[...p�b�5~Y�-��P��p�_��w�����w�����X�|���g��%gyN�&P��#��m�&#��Y���`=����dT)�p��d�,K��j�JcC�v0��Wy��� mT��UR�����f��T+ں!�(�Ӵ��lm�mS��J+�u�UZDB�b����z��%��(����op������5:[Q(��Z�m�Le�SY*!u]�\ph�C��K=DWR"8�v-��H�`�]˛����,�������x�9Ys�ܓ�cy�w�az��1;����܍Hz���c]A�Jy�Z=S �����;��?:.��]���_c�%2vN�و�[mkǛ&� �v�ߥhn)�/�S�	s�Q����@�S�ARL���S�Oߔv앻#�(wy��;���)ރ�{⇞����=����.�����y�I�Q}2	;�l���Ѐ�As��٤�o�ǽ������l떲���8D$��#�wz��[Oń��[2y|��x6�"�e9��f����,�!...��S��5�����<����<e��iZ�uJ�")&�t����w�ż�U9*�d��n8}�.��%/?���>|�j[S��K�bUb{S>Bp�(�F��v�by�����Ʉ:��֣�	g�3=?g��|��������V���M@���b�U��Wה��Q*>}uɳ�BV$�������������"��i�%3AH��5m���'��٧O�^�U��7~�o��wx��D=�G�%�i��d�է?�����Y�4�    IDATa�Z��//�˂�����S��mXm7�Ր$۴-mS�X,�뚸j8�j&�	n~�[��]~���/(�<"�ȃ��_٬X�|�G��?��?����!3�gO�nZZ��������9���d��L�:��)4�m�����n�x6�5�z���Lq턳��M��O�������J���?��+^��!lM��b�%��V[����{�ɍ!��S0��pu}�r�d�ڰ^V�@��8eP�$��P|�]�����_��f�l��g\�xJvr½bJt-�h똙$up�h���н�]�Q�ZOӴ8Q"��G�`��s����|e#�pE�+�	���Wcgo������}����٩�7��!4ٍg��%��#��Õ��1R�q����c��T�ػ���vc�{T�q������}�[���t�Cƺ[DW��I�#�[!e�S�	vJNqU��مR�����p�.�@�4"e֧r��a���^��xW���+�/�����T��`W/?��oǷ��G�`���!�E�]�#t�ָ+aO�k�aK^��9�͊G��9;{@usM�<�[G=�A��������dK��~ǅKW���w,�3$G�j�AX�����A�A  PZp��pgvܵ�\����É��̮���+3��	���5�P#4�i��YF�h	MG���d]`����)�5e��YJ�e���u��g�^l��u���^4��0������r����Z	�M >@����%e�\C1�p�;�e|r���hf1i4OH'#�R��w�����$I�(EY��8;g�Zl�(-(��:<e6UHb�L��+/eK[YZ/Hs���������S��1�bf���9/~��s��J�Sܻ���v��t8��֭H�ί��ox���\�W� �}��F��	~v�҆�y�|���mR)�:��.&4�������G��S�����9�?z�x4���W��k��IS�cH��Y
8�}�,U��C����8~�y�1�ME6;������/Y��OI�5��RA�#T�Z���eSsU��ʐ���h�m]dl۸�jI�j�r�Ã{d��YF�x89&}��d%0:�Ν��.�9���p�Yf�|�U5e]!t�����l�x\pxrLZ�X\]r(b�rkS�P��-)Fb4�,͸g|�?��?�s�����6�O������ڎ��A�Q*�	��QUkTV���P���RH�	R��������k��9���rh#/zE�-��>l{��/{_H�&��F�aoΛ���~i�x�[���P�0����-�0�m�z��j[A��U^�@������A��4�� ��Q?z���!l6��#�<�����^��W\�}�{��c������Qb���vH��.����!C��k��ii�qm�lǧ�!���o���x�>��kq�|�[�nw����>!D�t$zC�����m�L� ��㾽��5dENhVWKFiƭ�GH�8?{�T���-e���ÂJ�.kή.9�JR)I�&��ѤM�u��Q���ڎy[S������2ҖJ)cC��:��]/��B*Mb2FI��3�YJ"B�o;d�wH�C'9�ܑIM�^Dh4��P�UE<y�aLB&
�"vv�IJ��K��Q��hDs��M���dF���mC
>�L����}���G����5��iR���_�րV,ʊ�����~�ܺu��ш��8{��7o�x����^�ؖ�t��񌃣)�:
��Ф�@�X�T�?�%<��Z��L��8�]��1�crz������"1RUל�������!M@�͚�)����@`F#�ֳ�+�R�5T���Z�4���oKݵ�و�xJ��/����$]Ӣt �&�	E>F�1�\#}���;�	�j���/������	���������� щ�b����<�c#1y�j�B*��l�B#�atPp��!_��w\VK>98���:O(����%y����	�?R�~A�ZECz�E'�o�� ��*m�h��Xd�ї
Y�(���v�7����6aƷ�w�}2sB��Wq���)�ߠ֡ϼa��~P��З��0��'�o��8�������ݞ'Љ:�ygP;��ߧ��m�Om{��� Jw�;bC�҉��B��D��`6ǒ%b3�ᛘ�qC6�������s��o�����og�o�+�.\�?�����C_7�=���p���^�Pi{���s�Fp��Sd#rU���k<��{�)gWx�!|ߩv,�i>��Y�<uW���#�G*��y�L�f�!6?qm��ͪ���e��)%�)Y����5��#&�)��\��%�k���&! �e}y���L2"%L'�ɔ�9�k�u�1����΃{���D$�.+��c>�sqq���3���n��%�Ҥ��5-��U{t�!���jR'2��jn�f�b�S�bĪmhҜV�b�����y�x�s8+P:�Z,Y^�!(��-RNoݡ(2�h�LQhO��,�IBP��Y��qBSu`@u�ų�>�0Is�\'��/~���|�h��u��h���yQP��m�k*��iaP�<��*$'�d���	b���*�����9��f!HlC2��Bu���ylg��{�6)E�Q㴠[k|p���hڦ�0)Zڦ$ӊ�$46�ڀ!ZgcY���b�x\@pX���#F��6@��W�������锬��N&5��.GS���y>��c����ObK�����<��8k�{�Auy{R4��Z|0*A�H�-|���Ç�����c�Cv�������Ok�/�������ٸ���*�~���ΐ�������o%oǏb�rn���rl#$��.��y)v���=�Jz�̳�-nLr�:��G�Ҙ�"��]��(���|���oKI�D�����^��R���V	� 	�F�h�L�x+,���[]JA豪���_8�q��%"�ޭ�߆��D��>�Ș�t5Y�㻈>X� 5�� o���뙭i�|����M~��m%��o�M1y��bc��\k"&�X��'����H��o�����֬.K�m>bI��	VAJ2!ojU3���
C�2�ЬL�r}�hv����͋�����7tA`����bw��hL����5�d�����"�7ۢ�SV��h��C�F��[W,� �3��+N�{(���(�m+xr�>����3BZEW՘4ź�y�%#���=~�Yy��Pԋ�?<�+y�7���\�����5Nu(/IӜ�㔑��Oy�3�M��і%�:T��F#`u���.�Ԋ 
Lb��Ç
I�o2KItF�YT6�3
�3��h���N����j́�!���rx|��*8��C�����y�O�������1�<g~��mU���TU�l6���;�O�����������SJ�f�&:���0*ܕ2��$��!+��st�RjM���;JC�rQ�$
R�P��.X�"��).��\Rsb;f��J��a�'� �')F��c���ǡo�5���\E{uF��q�Ř�4�8�2�Z^�]5�u4]�A2fRL�J�`r���
�ɕ#�L�1��/y��S�b�o.�drFz�!˯^2j*��ۡM�s�G(�2)���e	.V�(yB����S����2h�(7u��*�k�p(��md�>�h_��Ͻ=�e(+�=+�s�-ټ�����^_��5IP��m� �Ï�S�?�;��y���M����Gqe ظ�$UX�#k��M�cC��t`@�=�=� b�,����y���:h�A����@����,��b3�>?#8�1<���,��
��랰����n���u����f]3~�X��O����F4�_\w��Y�pa.^1x��!a��|;u�!!�zOՔ$EF�Z
��u����*�u�)�P<�}V�M/۷���{����y����F'
ږ�,y��9��Md"s�"�霣i[�ԤE�h2"h�zU�'ׇTd�q�q�.�xl�Q�������ׯ.�<yQ0�2�Ƹ�dr�t2�0�q�,y&`�'�&��)I�T
�F:�4=��$�w3yJjr����� Z�Mg[%�lK$W/^�������)9���YZ�:OPn�A�4�'�%��@h�IA�',E �H~"�&�X�2�0&��ey�=2�G3��1F�,e]�i�-#��1�.Ԭז�jI�6h�zG�.!��ږ��Y�n�͘NOx��!���=W�ͻ��!&�	'Ǉq8=!i�\�ר�ùH*�Cbi���b��a\�p>�Js��A��i�g�}F�T\�y��՜�tF�����FcD�����fS��Q6bR�LJ��zB�:�L�B�Q/����46�qr�6i���!�^-,���r��C:'��zSJi�!���׶mo�JF��*>�e]�;A����W_���o��;yx�c�r����jF��s��B����H����}��`;�rO����l�ܶ=ݍ��CK���}y�>ž/'޷���u��������}���� ������u���<�&8{z%��m�M�d����7�]�jq������뺮睈┈0��TK���I����&/@G㰁�w!��Z˷�9���$���nN���]ohH!�J�4"�?ް�빮o$�s�����M�M÷Ef�F3_�1�����%*->8�ۙ��_����yI>4�M�I!6�l�Z}I��`�5��t����sx8#�g�痴e�8���4�o4!^B"󗔒v]�E����I�~���������)���j�H�QU�V+Rm�u�'�w8�4�^�Vd2�Lji�[��}HPBG�	�҂W%ѣY6E���p-��9�����w�fUr��s.�����_�~����1ҚB(��Tt�`#���3���! +r�{wɃg>������%(I��x;NN&��(���$!�s4��(.W��rӒ��e*�>G�,�s=��l[҄�ϟ3�u���!�'?�	����m[f�vdi��<�Ȳ��(��P~����l��R�qTli�4B�H��N��P;�2�$<|�?���Fi���K~��_�X�m���" �:��)GGGt�a��:� �ƴ૞�(�$"%�UUa��� ZI$f|ĝ;�����7}�;�-��_~��=RJ�E���x��%��c�阢(br\�P�)�4�#��C�^�?9"Ԟ\S����ҩ��N���J9�>ziRႠm[����j��]}s���o�ìۊ�CN���ǻ�ҷ	�i��m�`3�{��>#c�ڮ,
��W������u�mG���b����=����u�$��置�WQxE�՗����D��y��l��ఀ��`���ݔf]?4ז�5�sӾo����C����^������T�c����=�UI>��Ԋ��d�!��c�wY��q��A]7[���J�{�>�߽{=���C	�ش��i)�B2��p|z������3\�b:�D�s��Z���,�$�d��	i��q�$��dJ�QJ1��1�1�ȯ���m���$Inݾ���9)��׬�E�\��'�0i��u�0�b�H-bU�ǹ���Eg	f�#L�P�/�ߔ�:�@�H�+�zMU�x��%Ip��Ջ��b���Q�Ѵ]��&���C=��M�L���q�r��z����9U��	(�ٔMU#� K��$ޢmKu~FUW(!���6-��TJ����X�k1ư\���Oʧ��5w'�?�����}���m2ʙ�G\�zI��9a>g�t�h��>M�7b5>I�R�&&��'dYFk;r������{���/�x���){�kIp��t¸�.A�[�g���4J-AF��Tx4-:4� >1��!��SMÁ�ӓ;�������c~���QEq|�1��j��r�X ��3$i���7i���"qz�������0c��1���a6.��pA T$�q^R7-Mm�>��y�o9B ���Q�MW�r�{�D!Ħ�从q�y�a�o�}����Q��y�rX7c�&�m}�{�Q��:��ns=�gd�hu�b;��؄�c|w8d�$9ܯ�BOחd�k�$�����Cֽ��!Ě�}��GȞO�M���؇#�φ>����[nb���XV��$n�چ1��ŷ����{<ܛ�Y�r*���A�*r��3ڳ�o�#z!�~���Kڄ���~o}���s��oR��f�췡�W��i7ﲧ
`��<���/.1��ރ;dE���*[S��xBQh�	M�	�u��|ɱ���1k!����h&�	J).//�s|��p��ׯh//Apxx�d<&O��,ѸeMhB݀�"�� �ƻ(�����KE�ԅ�x�Ak�I�I�Rf���,�Z%�J�!%�K�O|�	YJ2�'5�Z�'6
c�!�H)MCoL�V+^�~��j�R�<-�M���ֻ(I�Z��5�Ʉq1A��c�k�ׯ�(��S�밾#t%��h��$�C�VdZ3�N�ۆ�<��_��|��ܾ}
����C�I���n�ӄɸ`6���u%���v$E�%A��q��]M/�m�.�C�$��*ڳ3n�cu�p||���9W�,�s�VYN�4��e[���	I����s8h�РS��`�E(M����y��9��y̓�O����𽏿����i]�֒��Cf���a�Z��PIL��L^�9<>b:���_R�%o�^����Ȃ�,�8Z���&�q<M�jyE�ed�<e�F�� PR�8�Ơt"�n�Mc{%�u,����濿�r�1��I�۾u����}�!�/��z�Į�a���j�����ro6�}@��J��e˗e�V3^���qa�߄6d�`6,�>"��j]d�"v�(/����^_�#Mm���K��;;(��,������77����4�a';|���[psӖͼb�!��a�&�k|�����h<A[	\T5�'w��������ů��5p�.�zH�K|h}����M!�w݋��~;�&®���\b�!�6��}����%Zk�N�8�}���s^-��F�&ы����!���5i6�0%�4/PAm��m���O��0;�������JJ�V��zQ�)�5f�*�zO�*&���]h��a���� Z_�dh����ݩ�Z��B��:���ض�r���C��c�_
VmK�u���	�#�'����	������4OX.����8�*�EAVL(����moP��K�9F*�"%ϋ���6�^�b��)��W5�J)�Jct
2�&��`Ҍ�jIq�S 2�FH	��������b�0�h!9���\�ueW1�9 ZFr��r��gz:��vtVQ:��k�=���$��s�4!�d:�������/�����X�1�)+��L]��Z��H�
�u$n鼣�,���'�r����[���iJ�����)������_�Fk��&���q�>��(IWV1YJDȽ�֑A�傤�ԩ�IO6�կ:�шP/`<AyC�Z�UKU�@�&)B��ʋw��m��.E��-oc3����mq��ؙ�[z��\2޵����\؜۶ݗ}ۊ~��W[ivʓv�}�5%$ND#�����{&Vٯ���~��Q?�ߗ>�/D�.��j���!"cf�\$�RCΓ���z� ���D���}��A�G3��{�)�l��Ds��ֆ��0�!�-�n���SxL�m�,V]˦��z����������ls������m=���Z�g�!��߇���^�M���OT,��(�QPj�e�����7o�+����d�[\��+�k�:G�y����Y���Aд�oc�#��C�<���	�y��!�''��%uY�Z-��2R�:ҧ*E�q�Ҟ�X�n{!)�ab���2VQHI'T���!MD,�i�N�r�$�1FP�kV˒�9Nf����:�ItB��i�H�3r�IA���	2&쭗+�V!LB��#����/���z���|�x<"˲�Hr����)_�b���T�teM�	�iN1�D�А9��[|5��AQl⋓ɔ�G�4͙�g��3�T���kKڦ�UM4D|@���N�ѹ��u�r�0�:�R��,�:ZӍ�$� ��� MR�ܹC��^�1�U��ʖQkY_^!�E�v���~��Q[�u��v���e��0t�)V�    IDATԫ5��h�d�!Uܿ���?�=�חdY���C����rCۛ�4
4I��a,%
���ǣ��|����`t�˝���8�P5���������9�����P���eK��d���P�Ȁ�z�}����ؗG��o��/�C�3�n���Iᯓ�v�I�v�{k��y݉u�u�>��D:�e���7���uK)A�ػ�{�<�k�P��F�4/�m7e��=��@<tŋIG�eu7��0B\ȵ�K��_罭���mow{�a����1x�7��7B�������m���gehȳ�����0�b�3�m+�ok�nwt��t��}��
�ws"J�;!��HJk�Rt>f^I�7���hi0H.Ηd�C�|����e�!��d�����s$�1���^-���&c���[�o��	u����#l���cͼ�$I�d2�k[ڪ���_��F�pB2��&1S���#�g ��su��:G���b�ib�i)c��Ri�by������g��?|�yLȺZ��Ĭ*�UE������<Az����u�Q��v��#�����H'S~�٧ܽs;��W0�2�7x�Z ��-׸�"E ��{$ڶC�)eL$KS��tm�z1���������k�߿�l6�EHD���۷o3�3�����(MU�8"ݩ2H��@x�4�͂P(m	�c�ǫ�\w��\]]��)�����<R
��:�֜���&��\��$�X���]�)E�e�����:I�2E�$h��|K״4~����ׯh�g6s<;@	&�)�����UUqpp��Zg�	���$f6�ͳ�v�`2��e)��
�%x�G�#F?%9:�6L�9msN��V�[�<1d�$ֶ�����rd��]���~��m���m�s�����W�h�m9�/���X�[sm>�O &v��m�'7I������)�gI��c�և���W���w���R��2`���F���"��������ִ(0I�k�Ϋ]�bk��,A�^ J�V=�gd��(@�MK[D��4fM7.�[G2x|!�B��.��(��@�)��8�1Б��x��Z�!�IA�����Nb�G�\��0�����,Z��w�S�$0Bc����B DB۶[FI�F/r+� v_!^+Z�]kl��β�~!�xݦ\do��M��6�2
����8��},8!h)���^����b��ܯ�=G$��~�CNO)Nf\5�,�t������> �j��s�x޼�w�w�K��EP���u��]�$ϰ�%Uǔz���(�2�w}p���1�q��%xM�& s��c��!�c�ҏ��y�ےW�n���=v
�m;rmh뎟��/���:�^Y
��ghj�j�x|ux��L>"	]t�Z��Y+�?��� ��Oh��5��$��ۏ����ڲ����!��m./ϙLcރJh_�3�,���_}MB d��T�`B�sy:�x��7�ɉ�4^�9�"Q�D�~}ƃ���IA Y��x�2�I�D(�����bI9:��j�v�T�^�!:M�@۴\6�j��A�L�N��\�q8��zh=W)AA�6t��r��cmK:�`���>C/���m�]��%��]B-A{����G8_/��HFb"X5А��V[���c����_��r~�r5'�!�c���8g�'�U���B�UK�Z�M'�㴘R��r���:{�ů����`2;��	֋ i2�1+?�$��������"K/�B�ɐ ��?�=[��1�x�����>gc�H��m>��1~o+�M�����R*6��↡z4W���y7,��ʷU�Q!��+N%�n�	�Z�z)�6�BFpA���B�Q��X�HLA>!�������F����$:�x��#1)�� 2">4��b�c��(�/�����$:��8,JG���asѷ.�N����O�u���v���D�Ǹ�R
#�xZ���mI���A!���m,�0���Kѽ{��Y�nV�)CS��c'aF�y�9	\/]2�����:�"����&Cx�&T�m+�l#�J$R��k0�/QrB�ކF��z(K�T %p���o�Z\1��ǁR�,����ގ����g���P\M�g~!���$d:B�*OhR#1�̕#��z9gu���49���xF�Kj�^�E26$I4�.�5+������#�޼�7��s���!�xʓ�:��ǯ�����ł�����������5a�"xK���o��$JEjR�q5�p�j���3\:e�r΃���+8�*>��'�V���H����)�k��13	�{�U�AQ���Ղ"�qp�@�+P*Aj�&r�+��FaRE��dF�r䣂��QG��,K�D�cE�J"����D�>����	��[$J��1Z��{�+�2��88>�d�`�R�rYKD�h=̒C�O�y-�<�j�S�S$6%t������ф����<��N�Zb�L�@'\��N�L9=:F����\�v$��0s��;"���f|�A1�|JZVh!18�*�/i����'��D�ljF�";:�r�ڣ���*\�c�t��@�7)�?EҾ/D����GA��<�Aan��.�5�e��v��M2x�q�rm��{��l˳�a�����.�PR@耔*"!v'���=�LD�n�j�T����N@gZk\���r��|�]���:�,Ù��\��[b����O��q�f��V��(�6�O;(�
��'$�>o����R\g�{�6 D�9�닼��/\��w�Vl�&(��u�;�J~���m�L�P�����Kn�e\_�w��c0.�w�� �*{��o6���1��	� E�������F�y�%�Qk)il����ӯ��uh)���T%�]����˗�&9�zI��/�8s��>hC:@x�Q}WD��<m]"���.�\�xF��K+Ń�O������q��Y�� ��l�H��>��,�
���Z���3�7g<��JiB�7�g|�������o��Y�H�C�����5�o^��N���D$S�����Z:�w\^]��W_r�J���f���g���$���	E��@��;��*������J�p���/�KD8<Nx��P_u���[P� ��I�h���M4�Y�ݿǽ���]�Z���^�)�y\�b�.6-�,�|��/H�	�(�:.��q3xt��d9��ʁ��5���TٽC�q2��� t. �ݗV�Q��h�I<��_G����r��8�b]@�)F	�b�2)�Y�$� �傧/�~�fqx����;p�OT�>f����Ay���_���K�7g<:fr|D]$X�b�x�Gwi�a��S^]�'Sm8��b9_E�o����>�
l��=Y7�m������a�����C����{[ކ+���m��_>���5���6�\�A)hi�\����=Q�.��l\�>�iv����%b�E�	�o]�������N��<8�/�#D�s��CBƄ� w�C�o�]rw}�Ǽ�ɷ�����>{{(�=\o�ݹ��-���`��oj42����=��x[e_��|dV�6^��F�vH�x˰�Y��/˶A�������ێ1�ܶ1�>�����⎽轈IzC=�(���漫�-�{C(J��`�d\5U����g<���mp�X2��*�x��MB�h-)˒�e��r�V	��IV��m*ʫ�ؓ]+$1�C+u]R��;Fi��r�.k�r��?�1��c~������S�S��	!����w�S�g�x����
S@Y̊)6�S��ri�
d��H�� �h*T2�����������#����J�X7�F{f�B�R/+.__p�:���oh..������!DB�4M	A�G)M6*(�1�;�X:7���>��	���m��C�"�B���&�9Y2��k��Ƶ\�yC+5�IQ���V�,�� 2f�7MË�8�KLș�?J1�	����IB�Ev��M���"(^X�\�eN�Y�6EH��r�ղ�2c�ke���(�X��Q�9�r���U1��ŏ���gt�>¸(�E�
��`��s�^a�*Aw�juA�����_���k��.m���6H!�������Z�Le��Ws�5���[��O�Y�>�NӇ����Fҝ��kdo[�2`[�_�A���<��6*	���2���{�2&��A�D�Im]���-�8*�Xn3�=B�I���bXV���P�o��P4����s���s�<�*&n��qЛR��⾨�Z����]���ch7��{�����~l
��2�ݲ��������>�\��|�����޷�Z6�l=�C�ǘT�	B��9i����.�k������U������!��o�_+�}s?>��x����$z�Ѫ�C�����r+��J≙�^t()1Jcm�RO@'�b<�K��Ҡg#~�=���#:JZ
��P�"���,��eUR�5A
NO�T��+tخ�[.��CH�!�� 
!�&.J��Ʈ-���j���gT]ë�/�{�_K���tB^��U����tM���lY]\2^���#1���=�k��KKp6z���,?����c����p�/?�F"��D*TPdF#�buuI�\��W�W�늯���,�,���m�� H0$��N�&-��bmZ���������b<���Ճ��u��DH�x�x�ik�m�ǚn�P�F�ۆ��JHo�{AH�,I)d�/r��|���ܻs$te�CJ����A"B��CIhR���[Z!b����Β����8���5��Qׁ���== {�1w~Ř���r��jR��M@A�Z���+�<}���g̿�=����W/�0�4�9�����/��ٿ�56�;�%�w�W�I��v��Hڲ��+��;���o���˙�Go��~8s8�FF������S�?<\��#�QYú�v�nR�Q6��	Bzֺ��,���$*x���<%D�'�T�8$�$
b�F��
ѷڎK�Gd��7o��PK?���g�����O��=P����!*�l���(b��З���^/�9G��Dl����>n�[oǠ�%��gȜ�6��񶡯mE+y��4K�1��d�h���e���7s�]$b[y��܇����7����>6�^ ��n��sܰM3�"6B��H\�!�@IA��]��<���u��}��\b�g������equ�o8��3�W�y�U�d<��~�gT�W|A��X����J��1Hs����LF�3-9g��}��g_r7�|z��k��5YH&9��Ԧc�l#����V���[_aۊq�EOZ��;�+vT�#�F"�B����������G?��Lh�uM�z�UU�|�~���!��
�>��]��~��Q��\�$:h�M��Y,iu�5T��;�DRpt���Zk� I�(��d:��Mf��.�㜲}�W
JU[ruu��i�o�6�]pU�^.i����l���f|�/���d�] -Ftx�շ�EƊ!$h�+�0̲��>yW˘��@�%A������W�&��0��g?���T��`�FB���i-	��4̯.隆�|���9m�p"c��,�9�uˤ�1���(�KV�^�t�%ڃ��H������ڣ�����^.�w���:&�N�f�7��������}�>7)q����`�����Hg[��@�����0�ӈ߄�"v;�:b���bֻ}�9z��9�-b�!�hG��E�#�X>K�9L�]�%�b�0��b�~n�)ۊ��q���ܞHY����AV��������p۪���� ׍߅��<@��Ћs��b��7)��I�9�'�_|��Aoy�.�&��&w3���oo��V�ֱ!K�tΡd,�X�VTU�v~�BD���ʆw@����a���f����/�ݚo i`s�����\�>��"]�M�E��;���1}�uZ��46��%b[R!J*L�m-�ƫ@W��������3��9�B�Xpvy�N3&E�����I�U�z:�ʯi�|ó��j���22�]Y����BNF}�d�)���l%$!8D��z�9wR����t����$���P�	��j�(W��c�n�$�i[b}��&!�	ע~Ou.%^x��zq�ٯ��'�IY��_��˧�pUGf<�rAu�[��I���P)�)��V_Isy�)��9&��M�ID[���Q2���&>��g4�g�_"ˊz�R��qԈ��bEY�H�0;>���]�ƅ��Wg��7���
�z�"�@����"&P���tMK�e$t�U���/�� �u���b}�d�^���L�(�r�(7L2Iv:����+LU!��6�ѥ�gw>�]���*v-���q*He������Y��ʒ������[�y���tm�J3yx��G�G��_S��y1b:9@%� �ф���Y+Ȕbv4�]W����i{�I��<�[+"����gf�}yHI�E�K�ӂ�����l=0$A"��_��I�DQ<����twUfF��Ê�Yݛ�scvWUf�eEĺ_)I����������lm)��l���5��.�-�ն�]��|�E;i��N���^ͻ��јJ�m���j�EBX�����q�㠨�Z�N�ι�̈e�f��̗d	sZZ���=���"m��]� 7F3(��y5������3��Kf�N)@�/�r��W��	13kq�%�2uJ��k7`�R���8oCA��HsS�������i���w�#I;j��q�)���o��_��wk]�W��$jި��V�����۾)i��2v��O��	7��$I�{�Ȃ�Ւ���D�����0����x������wࠎ~��fN����;��s\�������D����*�����7r��02#L�eL�O;�m�rf=E���'�?���?�W�x�G\�Y�'��cY4� K���7�w8O���gx	�cN���x7b�ϕ������� ,������?���g���CD0}|�џ������9?��8 ,�9�1޿Eb�?��-dN��x�#E��*{<���"�A 
�y�=�̈��ӟ���?��ӟ����'\�y��9 ���������k��޿���Aw�8���/0���8�`�.ϏZ���c�4��FHN��٩#0"��?��7��~	�o~�3,��7O�1aI7�q<8=�Ϗ����q�s.�r�4:�yz�0
�O3��� |�?���w��3�������>���8� I���#>�;�>=�-	�޽���=><}����_�~�[��w���i������ރO�?A�Rw8�pw-�$�WBߩ����N�iͤ���%���7�i�k���-��I�1\%HC�NWm�ў�f���K�=��L�@T��J�[�'5���eL� �V�t9oFJH�ih��.˘�w?7�Kq���G��쨽�)���CHO8����U_K�z�Ym^�]'�:�,@�:0@ `n@�* K fD$L�x��R�	S�wf*y�	g0�� ��(�	�$�s� �9ǵ;�4�$'@�֫��b6=0�5��s�C6s��U:8����Q���!��=A����&r�Jz�v|m!�k�!��2�eYmj{'A�Á�M�};@�L�u�(s�1.+Θ�a	2�>�5	�b��p�gZ�vLZ\��i���;�|�<��A!�sҜqHH��:���;i"�9��~ƴ���������4����?`81���Π%!� v�������Sē����p:b�#�9���]���!'���㟞��t�p�HS���CX�oO\R���4�����x>c�R��?�K	��~�-DwI@4kd�'KL���Oa�s�i9c	xx�����~��,�'~���Ņ���Y��F�8`>���՗��_�SD�fa<�z�+��sHKB�ɗx�����Y"�G<?���ޛ<x�7�5^��x��������8L_�������q�`�    IDATDhiV7b`�DSڊ``��2���$ͧ�\p7:�w�8c�܇� ������-N!!�n�Ñ��#Nw���3����������$|���a1d/|>��b�3�$|L	?�iuO�K���xT�9�-M8,���c:�śOO`D��xϸ����������t�������[�+u����֒=��P�&.W�Y;���/d��9薄�F$�I]��i�T�ݴD���ύ��c>���\�j:��L#IE��v��89,�e��s 7d�z�Ï�4��Ai!{�c�PN�j�#��8<��K1K'��3:����iZ X�v	&��\�1%$h� �c���hIHf �� ~��19uQ+� K뒈����:��^`L��B��0<��gl����e��d�!sU�M)�(l�v�	�]ac�^ٙP����J����bT�8c]�ɤ�-i{���߷��&�)0�c�~�40[��.�q�����*���NE�^����= ��y���=��?�ܽ��4�\"����r��(�u�dH�i�����#.���<����;\>}���.>��{N�� �0�.x���3��#�����✃�pw| �d	2C�X����8@�#���g�ő2��<�/���0�0�>�X�`qG��a�'�55�HJ�S�)8�$�!H΃�4!�l���z5h��N1��3<{0�a�cF�' &�������gE��I0x��#�5ϐ`	#jH'� �D|��{���㋿�| .@ѿw��>��go�$a�	�'xbܟ�d$M"X��)@b��y��a��S�gwGE��7�H���HQ��e�8L#<? qD�K��O.��x���(#�|����x Ma�T��g�lr����Y����;8:"��^0a�	�c�������Ai�u蜢��)���>-�y�u�R����\�&��~�*̌��qǖ�U����E���ϫ�6-�d:`�/�
�[�PՄ�˾����I,TLF��1��	�&F��r

3dJ+�8nјg�A �b �����z�� $!�0@YIMPb�@�io�����sNP7>���}VگC��y�W_,²═�P�j���U�-2�r��T�Wpm��-��0��Ll%������*�Ԡe֙���6P�#���qa�SZ�p7�<��xA�$��w�>~���&.��)��1_&�I9��4��"�����w�0,���	�_�>��5�޿�7q�#�?j(V���#������t��y����X4T0-bvF��`�\ 1�#$�8�p9k��{���oqa���A3qyvHN�����x����� ~���&I���5]!x^���Q�R^JP�R�|8�oޜ��Q�����f�0R��#c�>.	��3\x�Ek�NC�8��0��P��zG,H���y���	�� 8?�qw<�SX���>�/X�q�h��� �Ys�3g�d*Z5?�C��,$,DX&ͯt.�Y0���8_f�%�$=~BDB�DD�x
�}�xN��3bx�p������J��|���>̇D��)��Ì�̘p�0���j9jFQC�j�$�М��b����j}�&�k"c*��\[��ιή��X��U�������{�3�KW��K_� �������c�ڄr�{D�!R���#�9����le�}�V����(}��m������%P���R3���^�� e6&{H�3s.,����aU8�WB�۷��Ò8bH#U�Pi�6Χ�"��|�D�2�7��櫍׎��`���r����HW�����F��گ�{ێI���o�ֵw@�X��ŞwW5�2G�R�$��<�,)j��x8|�/�������hiN�y� ��b�7ˇLhU�9 �K֜Di���9�xAJ.��B�����1\��c ��7~�������s5&K���A�2/i��zYT���AD�.��@�	��gSB�פB\� :��[�w����7p'��˥�}n�"�eA��r]��c�c D��#$A �}"|�뿎�8""�NX(��p�w��⯽{ ŀ��3ށ�V�\.�������"��1�~y��|�a�4�����w������O�����	�S�H���[x|��iZ@�L�l~���劈������3�qħ�!�8�N��7�b��p��_��8|��  �Gw���	o�#���� O�L�0��r���/0�s�pv>��Is��/�<ň���iSU�#�8��GXH@�^4�_�,��N\�۪�۳�2�A�_��W��$��}���3�l1 Tx%�>HY�k��U���2��"ش�7r����	ժ6YVE�PyĴ^Z��(f�%M,V��\��_��Qq��n�c�κ�5�n�FW���IɌ�7�w�!��Ad7�H�	Q8���d))f��Aĥ�}J14S����T-Յ�q���s#68_?s�'����_���K�&��s_UK���'�n�v��*��Gw	�e��#�a Q&���o 
!�wmo�[�n��L��?S���J��y��������S�8vx��i���%V�ȌA%����}��d�D�"��#�p8`�G9���q��O���>;y�ww �~	���|(c�8b�8%����)%8O �/¤y��q3���#�b,)���9������{?���BH'�{�r�yݗeAX4<Q���T	 ���{,1�H���	���������]���;ڇ �0�!�� �bv ���PB��R(ɟ\`i�8��o���'�1�9j5@����?��?��p�D<�q�f�x�p8 .$�D�iA��1��{�^ɉ���3�e��t��p@�Q��1><����G�@ q<@x���~���M��H���7x��q����1���A��B�tƒ��XLV�j����_��/�B���Q��R�C�@�!�����"�"��'坥_�9Xd�wW��j|)��{�����8�����;g�ջ�@!%t1������W�%9�H��آwL3R5�V���J8�d�hW�L������57KբR_Kc	)]�:��e[zu��R���l�f�5�Ħ3�8TG�ZuҪ�׋U)Z�A����WV�|�}e6pC�l���!Q�m��J<��{V'�F�o��~×�H�Z�J�\k�J�G�G��_��wZn�J5���;�I?�0����~�����o�M|�i����c�9�2�_E�VM��0�
��\f�n��b�?�8&����8���$��4��9� V;����D9G 	�1�˄�P���|�5�����x��=���k��woqd-Y�< �3FfĴ`�1����I& �(:~����u�i=�� %#�r ��N'Lˌ���˄�<iXZX���'���p�w9�w F�ڡĚ&�	C>���X;E�2<\�\��̔f�֯�i�='�8#� Y�����pt-W�a�?��I�٦�3�`�� ���a�����q7�7��!x�{�� �����sZ��㞀a�0f��흞_�z��)�K�jSi!�O�7�p�,x��"�c���.%p.nb��$��$�p#U��{޼�;Z֟�V�����9�
�������}ۮ搫��]�����o��綮�1آ���<�����ibr���\m�dH}3\�d�Z�R}ۻ��iVW�CB��ojO$㍬y���>�A$��n�Z�+���YK�B*�,�}�Y���#CJ-dfn��׶-QkMkTj���K���R�r>��a����4�]P��[l�q�__��)�#��z�8s����V4����NvP{M@�����k�DQ$��AmET r�ԶZB��8�������_�����,�p'���' Ha �SQr��I�0e8�	�8*r)��t|�D�8p!A"p�D"�� sN|���0�!K	�!o���3������e�hy����b�|�����{�C"D8�#FD�(x;j.��7""b^���a��+D�j���!���E�B�~f�?�#�3fGHiƈ�Ӊ � vS�G��#�( �H���h�����i���0�	�D���9�y��0F/1!,3N<`$ ������XsM$�H ��/�!�v�` ���a>gs��w�)������91с'���B��A�o0��g͎�� ��t $��E���k�$�pT��Xv�3A�g$��wpiFHO�:p�=\�`����!��ֺ��< ���Z�`�n��Y滭��֜�����o\[c��5�t�v�6��hoi�9��WB���5sa~!�t�c$�����*�S�
{�9y��B�63{�����E�Иo3SVF& ��*^��_#R	� k
�g^���1B��ږy�lR���R�z��gh] M���"���w��I��r{H�Epz�^&�WDX����xW| Ri#%e_t���s�)l�X�!���Mء�R��V3����������^RwY�!������զn�(pl���m� ��ob9��^?cܖ���������O~�ʂww���Og�O�hl��A��$�%'��t�UER6���p�D�p�����ǀ)��W����0b�k7z�-Q��P9�v�����ԓ��g|��=bZ���#��?��9����a�>xC�	�OF?������	A<������ו�J�<5�*jIi�!<�� J���x�;�0�wAp-l4�Q��,X��K����z�� ό�g�g^Wa�#>L����#��OO�@1�Q��5���p�q�a8��;\VS[?�����|? ��o�q��yƃA�D`�9^ ��9��~����IB��8#��1Og�Q�M@4����Dn�Y>]h�Q���`6�d�"'���������ǿ�{@�@�LR��nђ1�v��؎n��W�g�Mś�� rMo]/᭾o�_��K*�7#u�����䃴;j��D��HylY�`3l��(�ˏ9�L��	̔����YFJ1��6�LL_k`}v*�=�)��A)3#��)Ja��ˎ?��a�!R%~]܀�|�\�euc$0i�h����\��b*�[s ������y�TH3F ��!|@
�q�w���Sop��F1��I�\��:\/�f�X�9��)"I $��")�%?�r
ږs�$����j~ƅ��x�nQ�)�u��۸�ҎC����E��Q�� [�-�M�,QՖ��0�}f����rZcfh�W-������|z��陰����$Eu|��5�44�,�rݞ�y�1C@�!x�sX� �>�x(s"�:��$���3�M%��?��N��W��go0=?��O
?A.J�Dc�L7+��13�-�o58˜�Ú����y	 x�\
�p���m��t���uȒ�ؾ $Ԫ�����Hf�ؐ��Ybe��;,Q%u�=�9$� ��˂�B��9��3~u�x�>��f�����ph�nR��.dfD	ڧ��.���y� $�uO�E3g���8�y���ii�^����p8տ�T�c��q��c�ڳ2��8�/�,G���������ÿ�g�3��C @�<��pQ��)
�U��ӖY��'��}�[Y�6 4�C�R�t'9�{�����54mE���$0&]6�e��iR o��%1�����	'�oW&�6���b�|-�$���N�x{u��$���	�)���C��;@��hjmA��DBк�<��F��6u �UQ�I�L���B�A ���&B`e��%�=a�ꎫ�����}��s"�B<��DŦ�.x���5^Ir�qe`�"FJ�T7#�a��$�vfCH %���g�s���kmq@Äp�6�`�LغzUP�h}��k_��2Q[;�ݶ��%���k��+8����1���߾-�~Cn�f��K�T�L���V���!�3�s�h^琰��Q@(�"���t;Ĥ�����p�"��x*�&�Wr� �9=��s�I?����� �S.���M.e髅�jv�QI�0�V"9_r\�ռCZ�Br���o`VLbU�ί��y�j|)&B5h�L�pCYԁN�CX2��4Z�������=e��$�2�LlNK,�.�7��9��PP&��#��}.�	���Ã{����'�SO�����8G�шgfHK���sZ����!(���dE�%(2�B��q\���>G��,��BEJr�!�KY��w�h�Αp8��D���a�\�x;ϐ�P�Lp5|2��	��%�ר���W+o�����wKh��o}���K�-�F�u�`�,�o��!q9����Si����|�*�g;*x֚-F��?jL�[}y�9��)��%�=qi�ը"�T�w�R@�P� �B4�!d��4��Bݰ�1��iӍ
����b9�m��v��Y�v������b*{���@����i^�N>��s�����_�iR��oȫ#�/�}���y��[�)����Ś�DR�Az�V̀dv��)?� �����\H4�>s\ $�<���# ��bx�V��
A5-�=�kZ�&�3���̣:eZ�'@b�9�z�F�bO��Q^q@��Ț'.p`��\�BA�4!8�!Þ��,�ř���Q��Zå0O�sn�JXT�-<�us�_Զ�"�S�����G�o����ő��3=��x@r��:�Y���L��i�PR�ƨ�"?9Cg���(�I5n/`���Л� a�P^+��ܥJ��6ˮ� pxRU뜫$
0Bs7Lw�b{�3v#����".�!=1�zcOD�p���p������O�<��T�j����f/ `�P�_M� @�I��I���ā��>�aulkx������t�zԐJ�'	��t�1zf�T��%B[��k�`�[ KE9�PUm�:9����`V"���^�hr	MV�@����Z"����Eƍg�靺�[ꩭ{�C�=7ߑd.��C]�v�]�9D~�_~�=��E�/Kq�j���xw�VB���ܸ̇���~ccD:Dj�)E�٦2��H�*�uc:�Tǃ�;�|\�J�N��'l�OR����Tj��KcG��Q�*Xg�L�,(ڰ���tJ1_E��f @�<��Z��R&|ɘ�kC��T�ȹjH�A	�\���1��nad���s�xí$�!��#PZ0���S �4a F�O?�	bx���	�o/Z8. '8Re���%'�����H	�K�nQ���9fPPXIDJ�ĕ.�t�����Id���UƸ���HH�D�13�Z��9�f��c+
�'��}��VJ�>/]/I�mx�k��^�eBO?�"�r���Zl�?Be������+l
�"4���Z���p����EF ��6���4S�����4����i�.�Z׆����lC4�7� {�#�T�j��:6K��S���,\�k={>f������!�V����e��j�7��S�f;����9��>��+ ��s�C�x��5�Yeg^{��'�E{�s��)��2u�& �ĤU��k"\�l{C��F��ڣ�Ӱ�����-�<��*b �g5d�,�Ըn#$3̨���ٺ��SL(���'��%Rg�b� @q.�)����d����N�l:�$�X3 L����r�8���l�sv����H�:�v�4�f٧ X>����2���<~���<�D9duI�� ��&숨a��ƅ��L�
J�!;�Ңf
Q�fE��<2(�c�1ER�]��8�#L�џm%$�FP�F�i��4�TM	(D��VDr8��Z�g��7�h���*�;S{����~[���B�>}���r~_��ָ{&��{��[8�]�L�Yi�]��7�(�9Dj�눊I���/o�@�.pQ'6d?�W,� ���Ku�q��� !��1@�kr�_�Fs���5x    IDAT�8���Tg4�D��iI>�x(��H ��kg�������o\��T}���2��;=���pK ��e	`�������D��ժ��q��@7|9��vTb&�T$��!�,�F�H���$ i"q$G�vξ%ˌ(#�Q5�ˁr
��$߱���V?e�E��jNpy ��"�,9'm�H�MU�g�WJ �\�ф���'U��8�f���؛^��q~. vSB�Wn�v %�H�iQ6|2(��<:uh�.m��12D<�0;P���RD �&��A��9�X���qɪr3�^i5���MG]���dF�%���E��j�W�&�3�݁�GBŅ@k�8�t^���"��@59�P޻F
Q7M�}��ք�W�e}�_:�{����%�{8�}�׌��W���m�jx�m /|�6 ��+h�w�tM��g+�����zCu>[��>q��j���
5ھ&��^�m-C��I��'��R�]���*��,\]�J���+
&#x)��i1E�ޙ}Dm�		QD���E�*�(	H��HM����X4D������^���9�����n��&�\��;]N�|	�9��s���`�t}�Z��U�m3�ת������X2|Km�XL� Nӿ�'�;�����Cv'.3�I���
s��q�`�1��iF�¹�,+�1�*�&�I�4�xe�%�� �!��ڢMIZ$��2�\���&�����3�vO��}����{�,��By%�Hꉀ(��� �+g�l�@� q��(a<�ڒE�~ Y���%b��c��i �)"�F�d�:��٬�L��1u� ZF��2H��l�ET��hx Wy pf L]o̺'(#�0h�������e�I��Ĉ�|�j�;�F�AXI�7��^����J���}�0�_����J�߹z|�]�u����ȁ�F1�s�e��w���zC3j4e:�m�8A�4��p^'@3g�����楓-}J	LL�яW���'Z½B��ip�S�4����4}��;�č�3�`U"�II%8?ZdTJ6��4���D 	B�L�c_q��el��ݷ�ګ�Ѫ�,b!�<�NѸ��$"��{t�w'8",�F	����=�x���K\�K�e.l>��&��~C�!�K�$�=�;N��K{��TG\��/�|���X�w��XҲF&��F�旒��$ ��S��H�L_��TZN��Q��S����<��@Prl;Pv&������,hf��HMe.�L�3�L�D9����P?��m��wS�Em�G���� �T���!�0��cD
����%���xG�	���'N�K��\�r�s
c���K n�/�K	��	V� ��A`�%��LZ��l���^��$��=H΋�A�#fx�u<�h!$J#N4��N� ��c�,���#�{gvS��X�n�<�U7�g n�{�֙~���.��U�л[��f8�p�e?]�+\�~+�W���|W��+��-A�g��s�D]	n0V ���0 1���8Y���
1yD���}�� �8 ��9
QՀ�ޘZ�I�D�#(&��D���		3Z�R����S�Lu�� �W�v��:�0 �?F�J�"m�R�:iT�ysǸT)I8#��{�jv4[,�  '�Q�z|�-Q	�m���ڈ�E/%�[h��fm����"�	Tl�>3Vŉ/ŢY�%M��*KH����L���@����Y����ps�cM�z<B��eZ0����oచe"**ͷ�la���S]o���{!��|B��y՝��_&A�KS%�l"�o��LfyL�5��m8f���J�s�u�Ga0Jl0ҊL`�$��#�0�qY�<��h�8iA"DH�c��	2xܿ��{f��7p��#<{�G��a���$"�>��f�+�$A�w�+.՘����ȅiQ�y&29 k���`MÛQb�H�97f@��x)��x.kvZ0'�����H^��c�#0�mJ��#��fUhi~ܹ��Ê�#�2^)U�)�[ʛH]8jq��f�.l��A"��Y�v>D%ĸ7!�U�Ͷ	�\a�L�XZ�D"��f�y�-�H���IK�OXb���$A5�M+]�sZZ���M	D'�����(F '/1�'�iZf$��e��o;\�����C��J�U����j{bh��k�e�s��^Tb�֜S��k�wb�����%�#[	:��U��mmq��}��������Rvz��kg,�bi�@���k.֐2e.2�&�q�����uj�RI�
��\[��y����s��0��j���M��4;��`���	r1ǀ���Ln~8��?!F�9j����)X:�~?��+t9Jt3�]��vm����_���7��U��u�}4�����.[E/y(�+������hf��k��{�E+������랬�O[�k�GQ�+8�%�����7�T�V��Y�i^;.�?��S�^ڨ�ߒƍ��ڴ�?]������B�-�@X���+M���iH۷}ޢ+e}�^�\S֢����o�kFo�#�+���_kFU"��gk���m�ýkS�׉)�ȕeK2�H6�[�9��5�I,���сe]֯�d��������~��L�J�mۻbl:ΐp{�(U�`T�Lh�5���3���v��1,��'fo\?ۏ�x��P���9��n�`�}�>i��X�Yq ��K�Su\���Èӻ|��[�% ��%�kג�V G��^DU����௉�6�k%����}����${8o��&#P���9��ؚ��N��X��c�Kf�H�k����sLӄ���
�	?`ȹ��3P�Iq"��k����/��3�<Gk�[t���3:��(;{�Jf+���M�������5�����:fƎ�mٶi�;0}��=�l���7�o�[�o����#�z��>�h�Ιٺo����Z�����}u�}���bBnk�1�٘Yv��}&j5�ܕ1ƪ)�"�&K)��/���{U�DU	U��JͼT���^�_]��Vm�8n�-P對�����9�~��[��o�T�#B�S��}��.�H��ڻ.�� iU�X����,�عv�nu&�!����=���!�.'lR��.���[22"}'���È),��5}���<� <s�j���T\K �I��HsS"�L���H�[�ے8���uf�zM���N�*��c��P<���{��M����g�vA�q�b����epG<��p�,n��J���-6���I���F7�+�^�{�j��U�{C�w����:��Dޮv�Z�so��˵'���=<�
^=��q�Ӹ��~K�oѨ[���ku�2�жH�a��c� u� ��E�T������}Z��,�a��^e��x�WV"���mr[7�fR����Y�.g���ت0�ƒ���ڴ���I������BNˏ�ͭmC������{!\à<��ƍ��F�n|�G�v���Ԇ�m�1��OY��r.�^�=�ǭ�='9�DJA�`�4�Hyw���X��O�<������\�8g!F�G$�C@��6o�_���dV�%�C��
һ�^�s��ZPh_�aha�kr������s-��M����(#�w�R�
q�J�B�騱Z3=�빰�������N~(`Z�f��"x�w\�m�L��o�1=�0�彊����m��XkF���l���ګ85���Y�1ۻ��J;�wy���[=��
����������D��k���i}��͒����C��gk����3���d�\��Ld&�W�~�=3���H�93���n|�̶d����ѵ����,�;����֡��[�l�=B��U�j����7�B�
.�Ն�\�"JE86vf@R���p) ����y�ﶙ��݌!�p%"pu�k�oj����s�-���T/�~�)�˭�\M:0cń��x������*2���qIu���b�������ie��!���>�um!Z�K�kR�#0)�n�lKVq�0�5ξ�������Y�kgW�c����N�3�Ow8�'��ݟ=L��������V���|��Zn�����yl���%8l���w-�e�\��o��/3�~{��_߻��2���|K8�jk�^���=5k%�3�!���* ��}#��F��tQ�� EP!��rBd*ɚ4\t�J�{�Sܼ�K�&sl7g�6��[ m%ւ\VR�@P������Ԏ�SZvD�����Yy {�鶆G�t�j�Vۀnn1D=�Jcڿ�	�<����]&0�M68A�l��4�J�^:�����.�Je����	snzm����M��v�I��ͯ!�Z�^D���y $HԪ�K?$��lk��G;�-��w�f��koo�[�`�
DZ�Ɍ$����&{���7]I�2%/f����E��͞X�	�@��͗�`>Ϻ��c�V\�qu���S� ��$�J.���X��/�^q�>3��)�x'K�VҴ�@��$�Nx8���]�Α���B��FKS�\��=ؘ�`�/[{z/Eo?���--JO��ƱG����c��^Y	g9�={��$6����a��/F����&�+p�Գ�u�o�ؘWkVj/o�0S���"����x��z�#n�m>k�WC������oἊ�^C4d��t�k�܎�Vϴ�����ځ��AN��^s�h1�c-u&̡`%��dD2�K�ÔD08��ϱ�T��(n�@t��#P��;��Yѱ&�Ii��׽���̼��$�/L���	X"���!r��n��؟W��״�A*��5��UU�ۚ1����=ig���we�j
\4�b�ۏ�~:з��� 	J6K;���<���wP"-HC��,J-���OU�b�R&ژl�W~C+����������y��ڙV6֠�_��
��'|ݰ&�J�K��It�\aZ�i������oO���c^��n��N��oMh��o�έ���D^D�O�[��V�o�P��� *Ny��J�:|����Ll���� >��!�N^Koq�tPX8C����$ $H�;�:�3�h�A(�*QI�h&BHN�H�Ej�*�N���sv�
�����f9�8��@���c.��ݷ�/�k1bL��t��1�=k%ܔR��E��m�bXԣֱ֪��#:>���Vps������J
97�,y���fVϱ�N�vX��T�ܳDF���J-&{R���}~�!�I�c���5���Ro�� �)��t
 q8�˰< �2">����]��2��c��k�<5}�u�o���!m+�bɣ�܊0�k�BVpk%Z
�"9�	�5$��~�{��h	�(�����*i`�X=o���0R]�#�pp^c��oa�98�%&|��xxx���>~�-��EM^�Br'@
)���Z��ے�^ ?1fDeB\�KN#[�
f�)yxLP)�{�3�U��?��T5/J1)*Bc� ����~*�� �Kj[��E?���&�ϖY����9�;�}x�-}��Pqzśh�'��fk�WnK�-� �Ť���3КÖk)�h�Jr���@�}(�V�̕+�i�ҧ�12�jt�T�"@�\�<�Z�>iN��I�Dps�%E{���0���UPN�镝&��	-UN�8��y+����I9a]�:��� -0�r���Ό�K�mF6A��aG�[k���b�M)僢)o9%�H��n?��M���Z��!��o�+x�7<��A��a�^���֖�����4
OJr�gH�H\%!��f��TYې��Tí��]:�t���e�7�l\�TiE9Z�M %;��|�;8à��Z͌���H���- }"�kK�nc�{�C���4��Ͼ��-���Uٻ^�خ$���G�0 P�*i{*��4�QJ	�˲"�$]ͭ�C����o΀Fh\�<���Q�ֶ�Pc�W�,���2��_����T�a~"�KP%���U�/�g?�-�_3����	y^��`�����Z�M���9��[I�z�-fhFŗ`~�~�i�K�ę�������RI�tm��/�r}����_�6���նs�mb������̶G�K_l�Y�{N՞i�fwn!���*�bN��l��l���/7�Pm�6��"�1�-���Y �*�[֤�gտ���ڜ��|��"���ۂ��j����>��5�)"�Jv)	b�����W�^�U�긚�9p'����"��q��������Q&��	.�Ĺq�!�m�8����e^"����~N���%��00aI	a�!9���Y/���~Dd��e{ƊM1k%� d��\�0�D0���] �+%K�H]��1ݬ��z�De��cD+���k@r��m�-S���w�a��k�y�8�1�ڻ[�e���OsSo�/���pd&%=oL��*�����TA\_�䶰]��-ӳ	�/�̕D����F0�~�hg���A�I�e�DEz�#��gC~�� ���~^��IϿ�~���yi�zK@��b�� ��5Q�Y�z[i*6kQ���ML� 6��AH��%85�Q[}ֿyV�R�E��9޺ZI��L)���Z�Q�]I�1	�*I��o\-���=��}m35m;���i�CL���ja�w�m���{[���b��j]���F����WTO�'��N@����r�v�l��Ǚ(��
k�gu|������+/����\��=%�k�X���j�E��i�Ԥ��׼S~k�
3�A���Kc{�Y�%���.���_��%h޺�=\M��<Z[��W�>6��^�K���%�)e�jm��J9�]�U��:�'��Bx�:3a_�hm�+�$�}���ZB 2U����
���&�jŒz���<Cr�M}�nJ2߅X���TY��⻧כ:��L�����J"G�`�c�����"O�=<�]���YP��v��� ��g�	U�6k"��U����deo>I���kf�|Շ�1��x�5U�=8�}ӂLt��~Kԁ�_�Dv/����ڿ6q�u�kA����#ZU�k��KgB�f)��ێA�R�1�'���)�*�L�(����iu��7���Tr+��U���6����]m�r�ޞ$eJlo:<cN5g�,��;Y�C5x]�Aa�# 0��6Mvc���޵��^sV�p�����{�k}o<[��-��?��Po��u���_�4۳)�D�r]�[�L��@�i��u�dᦥ�6�9�����)%חoqv��D�� 5g���F�-������k����%!�]C�54'tAF ;ia�T�}K��z��ey�$��kM{h_��.��-�-G����~����Hin�<D$�
+�f��%c�s��t�_8P{�`f$!P.FR�H�����w����KL��<�ᜇD�������o+T���aj۳�[��g{��ڷW����n����-��~^=���"��	0�:#�EH\.����J�ք[5?�3�)��Q�r�"D�$�*	>[�$�b,ZkA�:�[s�}���*�u��n?o	@��仌�}��L}������1m��vn���ψ�ë~n"?
O^ӎ)>X��qB"���w�5M�=s�R��x�=�n��0)nT�B��3Y��+���,	@�W ��B�0���]Y^"�g�0U��G־������;q�[Ȳo���_b6Jj[�lKD��µ��>Za3Kcv��-�Ҿ�&��g�eLO��9/���k�pK��w�q�=����=ưxKfR����Ͼ���3��5R �� �DO���q��/-�鋱��[�|��陃~/���1s�ߥJ�FN�v�[��y��FK?�\6@�@Tc����(Tdc��\�?���Im���b��q�A�|2�Dj!R�V�\MA��5�SG(^�o�=��z������{�ݗ��-�ն�������2�ޔ�����1�=�mkL{���q~A 4_(&�L�y��4����h|�x�o��:�3vw^�߷�R��JK�A8f�sp�R˥��`l@���O�%��%�Ԇ�u}�=ΰ=���yYJĚX���{���ܶޫ�P����u@�H����-Z����`�^�h<�E �i��6�R�T�v?W�]V|A^�k�{}�b���c4%��    IDAT�.h��6ʣ�Mu8����$�?��?�����	"�y�x<���l�PC�{����B�/!��Hǯ���O��-�.�h��_�o��u��Kr\�f�c$aY�_�#x��M�<��ߛ�La³���c����V�Z��I��b�P4g��<��'v/]��&^���Dq﹭w�q�bF_�S�W�C��^l�}�q��{篟�1s[W�=C��-)��*E�i˄_�����K�(�w�T�%͌(��DTߘ��{�`���w	a	 ��|G\m]Q<� ��	vaz^@1�tdHr�%��\ɱ����r� ���S���ℑ5n4�.�ΐ9�!-�?�4�yPլ$�@.��xP��M) ���s���UPl���Zը�iG�3
�m�ў'+C�`��	���g���~����%�=�&� �N��2 �Sӧ��-�]#��`g�&i{&Y��y�����^�;��6��\�V�' W�:�jw�vMO�H ;���G}��U5�N���-DJD�60���������""%�=�p5'#�-#�"�{��g|x����;�C��=��k>��
9��S���cj+�;�����Ƹ�D�'�q���e濓�@1y�KOM����r�;}�WK�â��� f���oNT��F
	�����1��l�9�p�*�)�[���%7߭~K]ۍ�M����WKd�p�V"5b��,�!H�i`k�r�ߞ�ԄX-�^Q�qk�֖s���L�4��WpIR�uN�DU;T���z,��sq�e8Va�3�0#ffQK��bZ�l�*� %@ڿ�1�P]9x\N�cf�*�iH�z��6
�s?JU�AA��߃G���o1��I�V�RJR bj��f�N'��Pu�6�8�j7DĤ�
�N�t����}׍S�P���ڔ��q��y��F'{o���[�z����+N�m�guZ��im�51J�.�����&��Lq�����.�#�s�W�;�!sҨj��0`"�>U��-U�i�[	�Zտ���M�n��i4?6��'�0��'x̸��|�~��'��9k<�����%�i��<�k�(�� "r�w�>4iU�m��v?�G;���1m��&3~���I�&��:�m���v�r��=����]+uB�q�/18���?��D �Ľx����3��d��x	V-�(���p�m&;Id�⚑�z�վ�a'�4s^�ʗݍ1b�3��6�Ƭ8��` �b��Hиk�����X��afx��2�NtI�bF��<א����y�o���o��z�w����Y�>��j��z��hF��l�9�����s�-�i	}oϵ�����ת���6�V9�.����Zpoy>[���O���R�Ǿ��U����P��B�D�*5Z�=���#�mΆ[��a"��e�͂f;���/�����b'�$H� Aj!%��HQ6MJ�$R��c�g"&b�m^�>�3�'q����MK2EI\$��&�;�\\�w���>�*硶�:uN��X7���g��ʪʭ�2�2�U�Fwh�BO���֐ǲ�[�R� ���#>&5��e�\�%R�W�������aL��Ǆ��k�w� P~ϙf�����^�)[�׍Rua1�SN�gJ8C6�m��׫x8(�����<"�m#�ԯ��(��P��h@��3SL�&XEe7c�=*�xCȺ����=ٖg�>�"�7
�
��.��HO^�?ƀQ�)͚�F�L�Ơ�3@��e�9O�hD���
�x��aAk��Ʈ�3�����u[D�3T0
�(x���mr&6e�%j�1����̮$0C�����R�f�`J��lR"Y'�q��"�𻜸�`gD>&l��A�u��F�|��Cn1�*%魉s'�s/��TB2�����n���;,�����&@e� ��S�s�6��*΅��(i�Q��5��]�\���mCX��0W-�L���#Cޖ�[E�Ko��ǖݳ#L3%"*&���4�q�������'rL�y,��)_y�ȅ ��/�8�I�r�l��d%��T��%���~�1�)&��8��,���:�~�hbM�-���y���8΃j�|�6_e�����g�
gՠ�Pڪsq@d��(-ǿDΪN<\�3_�������j �Y$�j!��j�CK�@	�;� Xk`�Y{�x	�{P�!������(� �܄��|���?���n|����u�+�q4��2
�%d����BD k{�c�,�3��a<��瞏��C�Hg+֙鞈\ly��,��p���fkZ|�ݬ_��rAFX�|��  �0�X���� X
XM��ƙ�}�y�%>C)Q���W;�::9��t��ك�ܭ�}�Ӷ�;3��H&��Bayd=#���=+���3�<i�068{��&�H/��.�c�*�Xj�;���[�b"� K�vz$�*��a��7V���q!��w*)X��`�g9fDy��?��:�J^�����R��L�ż+?�|
}����̫����#l�*NZ�  B��i����EtIH$ @� �w�1l���:U�	��[|b���J���� ����fAe�p &_{f���⦷Lg�Z5��f�vٿA_
���=0  ޘ�袋���{��(h�q��CrE�:�av�i�Q|����ӐgЁD�%¿����W>""��$�p�=�s�;������L���eG:�֖:��t(�0��ָ~�4}ۏ����;O���mx��Z�Q(в�r.c8���ق��s�9i��� Q�vF:��Z���YBJِ$��-�8��טz���R� .>��]~����s7[Ƙ�d�G�
4����$Uzzc�e��7�'9�3��݉i��uȺ��ֽ�K:��z�¼�sb�I�`Od�钁D\!��6 j�\�.��V-�;��H#j%L�ˠg���d&�82	���e������Lk�f{'���7��J�4�=�g�!ʉ;�N/��P��aJYj��4��z�Ǥ�%�Nz�O����-�MM������賶b��
ls�⧵�LsDp���u�F�����c\@��b�D;)t��:��,�]��1�c��v*p�|B�2��̂Q>#	o1^D�Z�x폿���	|�?���>����V-vN���x�pD�6L ��'V9�w����-��f�������q$$\H��koJ�ZcI�����	}��!1��4��d�2& l�^�WS���~�]y������98�=n�/�-����P����{KQ߄��	'^�5"��ܗ���ڝ2E����;��$I��Y�I�u8����o�U�� ��`;��]m����K�tG�� n�0��Xk�i�X����]�!q��rl���R�n[2"$����ϗ���!�T��� �H��͗B���F0$���D�ҟMN��iĳׂ��Gw ���h�&4	��"4Ґ�K�7i�����W;\�� ���Q�u@8G�M�IQ�4CYd��Lk� �,n���x��~W�/\��bv�r��jp)N���f�)a;50֏)mH�#��$Pv/#�����zD��r~�1,y}, V�c�]�!_ӹ0�����ύ)
���Y�rJ��]��5�v<F�o%�낃��vk��l߽3Nz����Q>���1Z��@��yX7����i�^ܤȆ80�SIdG�"��WXə��]�wAKᎪKX�R%�8�IOh�	l�kJ;b� i���J.�N18(���Rm��������X@����mcZ�_y
�!@�4�0kZXk� �V��)��s\v��VXG��FH���R��&�gT5�&�of�ǈ���*�!�n��ո�jt!�80��Yk�2���� Z7 � ]���%f���Awr�Z��W�����	fD"�Jc�K�  ��+r�8F毤�d�ȳp��������Zk�V��N2P�C`��ȟ_j�Ov�1E-�g��	F�1`k���y�?7'b�r�����*�w闃�J�%X����ǿ����}�; ��ѮF��'3�M�<&,w���*�z��%O\3���J)�n��8s�� $d} �n�5m����~�����Qx��y��s�襣�%L��\����]�h�.؋�A0`�� b H�9����DGƚ�.�����p�
3ǭS�v=MU
��X��m\:T�4[�~��B+��a���Pn,xH�"�W�H&��,�䏩%�"�&�	��Ht;%;�<�G��������'>�:�Y�[�ԍb|�����P �`k�Ф4N!���2�4�kf����#1`Rq=6�k�Z�=f�f3�c�@0������cŬD��i�Ƨ����+�D��vg�w2Y���5P���\�Y�H��h�U
x
�X���yU�4q9���� S�e��PY�+�,b�їZEx�.{h��� �p�:�R=�m��[�����i|���{h�3caO��)�E����}t��K|�_.�\yT�����~J�)9���
�<K���1��M֋�^F���>#:�� �QO�T�9�*���%�����3K�Zƕ�7�����p��:*�^�'� �F���^k ?��uE ��N��h������+�3�tH�쉣��o�(k�\�y�;�V�`*Ic��7Q�L���B�8��ٲ�=iytrg�\-`ǚ�� �c�f8YZ�z���Y]E��(JTD��|)P�@
+�wI����Q6YZ�u���1�v��i=[��Q���4u77%�Jj��B`�^���4r����T6������ȡ�8��Փ�Gj��r4��B���&Kq!1�#"[΁���w�^2���.L���L�a�ëy*F�Oe����^�� �RB�<�u������H X��z�����i�,v��k��5v�wpp|��
������7��}�}����p���X1�p^]:���&��H�^���x�i/=�g�V΢�ﱢ([ԶhJ3^y]��BZ����~	�1{ ێ�֏�CBμ�$�3���]���3F�����π�����C"`�h+�^�2:!T�WY�Q��!T0o�7Pß4BX�٤�_��2����*�JXktF>��unO	��RSd���s���y�`�|l�u ��xf��Zhkp�<�j�����������1�d���oh�F3��)�I�=�|&�-�7+Xl3��Z5Ȭ;��H&��TJ�DY��q�}	�-�b�Nx��i�{��!��`C��)'lb��N#�$���葍�(-�Ԏ���a�q�|��|����HF/$�*'����1HF�\�X'��<z�SX j O�؍cn7�9ٙ=���t�Ƣ񺅱_�{~�Cx����q�}�>\��p��y�۹W
sF?�ܒ�Ax.0{yVڅ��hX/��^p!�xb�h(E���%�;	c�|�˒n3͚ݬq�~�C�6�%瘸�d�/,Z_�Ð�f��n���[��7��[\~�<v{AH���Z|���S
27I���f���B7��:{�r��_/�.Y��DuM��֔�@8�hwn;%�f(K
8�d��*նI��dQ�����+)�4��>��q��q4; Z4f�Y�¼�G�V.E�1��4���s���(&�R4&��1�|�=��i���>�PB�<��\��0����E�N��S"� ��t�u�b+8�-�V���Dhܞ��:��P<^G �|� Ō>�5p<F�s (��L���gyv7h���G��e�}�b˾�Ăm��U^�m�#���T_�6嵞z�5�sr�f;;�����GX���x���{\:s����5�j	�KP6��9H���t��X3gǽM�� �r�CQ
�)�)�۠�b�N1y�P���I��W�bd{���|a�Jo�rL0��vU�c�����x�ӟÂ4�7���y�;,pNWB"��W���f�wD�����*�����|���#WZ1�C@v�� RD�?$ĂHM:xå��
�J��)&��y?�r�j�St#�N��B9��pKa�f��$8�c"������~�M����<n�A|��O�§��
��E�V��Ŗ\)
����XE6���MQ������d�8�t�3	���*.,hxo��Z��`F�2�0QZ�9)��j4;ӄ���$}�%CZ&� Hކ�A� ���!Jizۣ�:����Ȑ��Q���6��B@�� As	������r<��i��KM*�'�SJ��[a1��ix�p������w����A?[�U�5���Y|��>z�
���'�^���bi4ñH��(�x/
~C�E !�y548/�2�Z��W
�\�E�g�j����t������s��$,C��(]?����`NNp�'�F�l���%��8h�$#]�'q_�;:N�w��{}�5Wz�v�%��Xes_2Y!gT�	�G�
�Z�А;f�@Y�(�nxGP5���ӀU��F{͙�����3��Ba���a�PPD0�s�[o��~/�܋G��8�-.|����Z`A��2�8f�A?�ⶥW�V��䭤���R�:��-���m"�r	��B~@
�I	R���A�$��{���~�
����7���z	�E�6ћ(�&a��c��v�5.�AjL��l̥�qȲ ���%�|��A�t��t�bL����U�&b���DwZK���D�$�p<���O�����@�D�����"�>�����\��Ghp}w����x�/�w�w܅���1��,>���
�o}�wv����v�)�I�OG��V��OB��=u��d��d�
�<�@8��9��� %�kZ���H��o"�e� 1W�������^ux��z�`m�,�`ae�5*FFt�A�0\�¹��	�+�����a�*�B�aL\�e<r9��(;LH�����/����>��ir �k5Mp 0`/���w�	�9�#��,B�{��gB��[���Y�����g�
:}�W=�N�_�����|�[88<�9é�l.�I�X�W�f[AI���sg�/�Զu�O�R��z?$q�G4a��e�&s?>�-cD.��<����u����Ξqm��A�1�d���1�c;X�am�7�Q��S3�h���K��d�)>��1�\�;/M�Zo����6rYgY��!Ө�:�Sj�)/z͗��OY佱~�f{�N�к��2n�yǻ��_��X�y?�� _�'~�_��W�-�D�x�-��fiM������5ň����BC.o9Y/���L�A�_|����`��ݗu��u�6	��l�gL��_����0�� �-A��k�0h݃�K���@��{C���c��N8�!��ד��q6��g1��J��ȈS%��X	�xKxB�r��*����)F4�@�R����aZc��>J�ٝร9���÷����k��h^�V���_q�5:��
]%�,�ZُT�$��f�R()�k�hoYwI�ܜ]ws5��Y(���Pj1:�9��T�PI�+�?<x���5-֪��t��iA��D^"����1891�;���a>W�ʢgw�-��OT����%A7��9�l�5�~r���r�zmѭ���6-�&L8��<K�@i��ź�Я�";̀1Bӎ�X\���XO�R��	��r+ར����K�иk�$<��q2(��@x���3���`;�s����#��vpp����ϡ98��y���_G��C0'G���7�����>�[��3���t3CC@�\�m[�w��.<�3i�h#<��f���Ι���ZE)����P���"�?���A�*��WZCA�c'P�RVak��טC4;@���0V��$����p  �I��r�ʨm��e�`n>֯q�R(r�<��U�F�+��3�-�n��)��D�S�cv����;5��LZ�0�H�����ZT����u1yջߒq�ր�[�`�1{�W^�ē<�au�Z�{���F��_f��˺�
���+�s���|��3�Z��]�G"r�	�B��Yx�ť����p��g�Ʃ{����>�3����/���e,���ͱC��h����~{z����"�᲼o�z��59�3�A�r    IDAT��1�)�=g��M���+ra���hƼ������-@�Xh��0Ъ�1��sJA������B�;	���T��a5��b,�BC ���*�LYX�����Ų't��&Ƣi�if��ܸ*"�ͥ�w:>�q�O��_� ְh�s����e�('�Rʻ���C	=!�f���,�N�S����>�Q#�{[&Ɓ�Q�T�l���D��R[�@ŹHܗ�Y�Ve)�p�_1��&�� �>��fѢ��Y�m4���!�g^����{>�O��{7n\~�����߿��w����5�����;>`�O�h��։^{M�;��4�7R�J����R�����#-|ɐ ;�q�<S��)�O>&��wK��ɲT{w
&.�fc��M2b�-�����ƙ��IP�)�ZM�-�[M�k��m���u�,-[�g����럻.#7�t��-���b�Lg�s���6���,�Nc_+���Oc�X�m��bvϽ���Ga�~/��|�s8��j`O:43X���I��'��H<�aw2�4��������^q΢I������	�L����������`BaiUE�~��p��iJ�)L��$�TJ����У��R8��ġ�p��ic`awL{CT���CA����yv�X��$F�I��+�rA�D\ٽ�@��}��I�%�&"�q��Xf ,z��4ԭ6�_� 6xq5ǹ�~o�����5X�\��×���������Yc�������hܶI�4�m�K���Y�j�+఑xŊ,�8I)�x L����G�hg��~*���@ (�s�x�9���T�P�u�ТPcc�Ʈm*9|�S�w�Q���l��9��G����h����=7�Y$�%�/c(�����R�륵��!�.r�D<����L�t@y6�VGdjD��#�����-�V���_��u�^�s�
�����O����r	�羃s{�P�����Y�6ñ_�# �K��sT
5᭦��1����՝���������$�y;+F�?��c�џ*�3"_��J� aD�v[9̪P�K�C��p��M�5<�`(�K�G)��*�%�)�e�Ц#2����R:�H؃K�Oj�)�郉TeM� 5ѐ�vB�P� �{\bw�����e��9$<�׮]��h�&oM���8x�q��C��so|#��w�
��;���?�Iܵ�Bwxi`YCi��l;+�ƻ�{��銵f��/0`*r\�+=����`v[3
�����x�ʱ�ʸ� 2	TF�Gj�o�dS��fJ��dN���X�����Q���%\ghE������Ȣ_}?Fߪh��LoL��ܱ�46!�B�$��X��`A�g�6����y����N;��"}�"�$i�&���y�$�,�,֝�-������O};�n���xv����8�2��G��K/|��Bi�~עYi�b����<�6�}PjJ~Q�)&?%t����|��H2ڭ`���.����^�q[������������5O^ q�!Y�򆔨R%�ޔ��0)��3h]��A�_)X���,%( 0zx)+j���l}V,By�+� �u�kT,�WR6zY�a.}Q��FD��D�M�~u����kK��d\����?�ν���q�:�\z��Ͽ��?����݅�4�NV�����e�P��hvv����z��r�D���V��bZz�'�/��gf��y��FU�E�٠�P������B����o`�9�����͖�e�e�I�l��+�*0�R�uU4!c,BZ�ic�]g`Þ�+(�-,*e�}�'jRx�Xr�؇E���i�˲�0�s�ܛJ��r���J��p,j���z��1Uﻪ6�?�ON@��	����z	�W�S�[`�.��,�=������{'f��)/�������sx����k �w�"�˃�bh���_��9-��5��á� {����|��T�g̹i���S�S3C"�&A����N:2[�t�Je}+�,M�ؒ��`HD:�հ��`]ٔY�1jx�;8z�c4R�pgb]��%�o��1��B�x)�&�6%�q�b
ן�D��o��7�(lӠ7X���h��<���~���c����KxU����'�?�(^5��t��Ŋ���g�������b���=1�<:v> �B���47��>��R��n������3�	<Ԗ�0��$��iC�R�4�9�|�I���c~S��R��j�g�p\\�P&|��l�2g�6j�i���7����b�:'#�ް��7ۗ(���Rc����%���IܖIm���m�q^zE{E��t��\�WR�BNPY����n�6|�5Xl�Jws9�k��@s���j`��߮`���o��o�H�����,ϜƝ��ih|���=�\��}&��Fn����E*g�7�'�\��!�/�֞���X���u3h�~��pwE�����%���-5
��9�"�E!ͥ�P������h���b$�"��� Q�/<�u88���˒vB V �P�����coMBF�7��\��hP~�1�m�`��0G^x&�Q��ȳ�yc���>8�H�G
�
��;��ټ�U68>���=��'ރN7��V��y�?�9�1 ��l� �����N;�V��v=V�lo�����G���~1�<V�dr콮A��"r��Գ4^+�O�!���:�r<���'8�nPB�xI�%��CP
���MR�Ĺ�sc��=�Qkϖst�� c ��3��F�JQd�cu%�W�*xR���%jIB��p��&��}�W/���J4Ɗ�%�{��Pߔ�}��>6��~���u�L����0����ʢ��~
 0kf`,�vk�VP�q۩Sx��3��G�f�:�~�ؿ�ո��?�K�_ą��3�{��\F0�0�����X��f��z,'̜)zSs\>+����i�3���NZ�d��r�Z�3$����,�yJ�TC����A7'���5^�L��B�.K\��H���ا@r ��$��^���	��P>ۏR*�pO�k\ �q�{ֆ�<�{��Z�3�Z�fd'��e�yX���b8�ѰFc�9i4M�þG�,~���Sg�/;��/�/��n�t=���]��
����8Y^�{�D��u��'�8��+/c�\���<ľ��35�"w^M'G�T��Q�ZGz)�q�+��L�c@A�Xv8!�����d��<ue(��06B	sx��'cL('FC�,��DH!<�r��Gd۶EӸ��}�c�^W	DI,�%?y@
U���~��.Ǆ"I�)SLh|�%A�~ׄ�a��}"�~�8%
2 [���'����0�n��f0W��e@��K�q�=gp����[��۸��pt����A���~{?�V��Y+s�>�籲�zHu��	Yʵ_{�ޮ�����0��:<-d�����U�$��Z�I���7[��U-z�@0Њ@��ѹ(�AH9������z�v�5
3�艁�w�b���	�(7`��EP�q��#.1q6p�(R�4�K��2ٱ���0 j|Z@�Mΐb-�r�!턐<66�;W��(�DP��T�)�}w��R/�/\�k�:�u�?�C�\��|�ֶ��W�z���z�����%�������1��q�?ƭ˗�������?��vk��
'�{��a��24Z� ��;��/0M����}GCp�I��X�fǫc�~�]8u�-8���8z����r�[_H�1	���]x��u&��i���P�W�ϰ��SK"���Lk�t繙��f'�+r֤0�2Ƹ�FB�2Z�>���@���0�J��p��OBR��pqM���S0mz'M�y�Ѣg�я�l�u�RCa����p�^��(�?�괞"#��;����&\��R(�a{' �ib��`�A9K��.�`��ƍ������&,�*Ͳb�ȿ	wA-Oy� ��Ě��źcX�0[h\��a���^��g����[�'o�Q,�]x��������˟����x�鱠=�=&����9����勩؏�΄�]!f��1jH�hB�n��L#�ٶm�,�7�X*�a������Pz�N�����&��`��)�5�x�}]:09G�����&ǃvǢ����W<e���)(��0N�s�F58���4l=P�ײn�aG��Yvg�ܞ��։|~Cդ��$�R
ݲs�aO�3�wD��!^/��%0_P��H����29g�,Y1id��R� 7I�cŽg<�.΅#'f��]�V�+w��Z�e��~�c��őjq�sx��:n{���5���!�������gt�V�p�w`k���`:ٿ���3s?��"�)��#�ҔDD��`���q�X���˃l�ְx�Jj3�����Y(-JCmO�ίf(�&�N��(�T'�d��XZ�OJnN�.�W	��&���ɍ�c���r��V���Ҹo��59��o���Oy�|.ocϕ�8�q����qa��4G~S��$@|���w0�,�}��9FO������������K_�]��9�z�<��_�g�?�+�~�v
��f�zt���0�͡צ�k�-�|8D~�K2�R��xa�5<��by�CP�Bʹ�$�M��	���x9z��$�!mp8o�J�X�P���czF�������0��VT]�a,T�܌]��@1�鞓hy`�w=�� ��݋ȑ���m��U	C�^m��ݫ~ԇ�E�h��W1��B!r��EH��
��Azg{x�C��[��a����=�g��c�ݸ�n�<YC��lt֒�_�����,!�E;� �PP�a�N�c���%/^�Z��{JZ0�8�f�`�t&��|���iЩ�|��8|R{5��v��Bw%-M�5ӭ�.�<ӫ=?%H���=?�fN����d�Sm�ڝj
�1Xkc_FE,I����`��x�HN�a�C[N��`@:R��H�7�鿄G���1E�Xw"F|3��J������?�����cy�x�d��7ԙ9ԩ��^j���S�Z�U
l��Y��Zc�U�Z8��L�_�8�+��J�����2�[ۂ֍�?,=�Xs�@���̇����38K��� �RhT��1z�06(Ƙ�R�ȁj4mn(F�r�$;'�VN ��tyhmp�o;��q�ҧ����m�
{uT�X��\>s.aa wsrѓ.P���ø�����Žm����������5��� ��X�������)N��n�x&������F"D�劙������{���<��0t� ��1����v9F��B��d&/�Űn�^��C��f����vI�б>W�ls�>C����E�"��N#��Dzw��^��������M��6eL��b�Su���n������}�mLBc+c.�0ȶXy�(��V��2����L��U=x�c��p��y���'��=8���x�]�]Y�pt��羅28�cu�}Z`�U֫r-�i���b^�9�)��|����)H�����vN�d�����Z:�ϴn�֟�A�Պ ۃY�@Ù�ÑXe�����"�z�"��?/��C5���&������g
��A�ɛl����v� �9��~���'���#8�c�����b�7		,�f/��������Ie8�G*@7X�����x��������)���ʧ�_��A-/c�j-�3��Y��V�]�ݝ�.ߧ%�7�X>FaR;k��Zh��6M�5�6A�����c�G����D�����4eP%�ȧp�ד�����!b?���|��B��0�L6Nl�B��6[��>����P24	�+)c�x!ڶlSϘP!}&d}c�T�ٗ�J��@J�p���u�h�1�����7��k'�B�.ɵ�p��:n|�S88s����oĽ?�_���?Y�.}u u��*P���m[�Ot??����)9��Ƴ�6g��z�wh�f�w�&����@����Ι��.��-93Ѯ�B��ab].6X�(�tn�1`,��
�bؾx���� ��렔F�= �/�4��~bi/�]}�v�Y�7.�r(k�:�=L���e7h�C�> �� ��1h��0������gJ�٤I���)c�~��=0���<�����>�۰�z�/�7|���K���v��VƢ��N�>9�\5�=�Lð�+Z�V躵[�V�����K��Mg�GY�APM�3	��ys�P��ZCNTKb掱x"�i ���k�l��m��̇�NwMJߵ�H+�w�a_�^�c	��כ��x��)�Ķ֨1�5V��Z��d�m���T��m_J�l�k���)��M8�f�Md.i��������k��?_獙��ڢ�9LG�ewZ�O�'��N����ƙ��}�|/��t	Gy{����3��j�p��:��1��ʴi|(�1_'RY�4okk��L���'���7p��鏁gs�T�%�s���Ki/��vސ���ѝ%�,î-l�;�E�6� ��_�}�	%��ݓ�Cg�G���0�&9RJ)k �D4pE�K
$��j��f����0�#g��5�ZM0�R��`��t����3w���[���y�k�o��_�`}��|��
��m3��;h����Q���ĺS��n�FO���'���`0���w4)X0���ǀ�,t?m��E>W/�`&���]w��~B𪐩xâ�'4ґ��
'���R�'�1��yY�ڽ�wƴ����R#f5x���P8�_3�V�CP**cǄõ��m�W�qDq|9=7�NwƽiAj���Q+�Ϸ�e�^/�׌;j	�����?ǋ��8p�2���x���ނ�4�jm�f�(�1�+q'��W��e=ec��r|���uCZ������ɩ�cs��&�]�ORX�'��Ƕ�����M�Sk�i��naTM��K	�'}) ���}��+�c`��x��Z��� ai�����d���#9$D��#7E:b�M��_�`�d�Q��j������n���?MNP
���1|0V0��'އ��gq�'/����it��A�-q�va�\J�f@��O�y��ط��Z��V�(��8��vǤ9�@�'x[p���%�1lљ�r��ehk��K�3���%0۴���k�K�Hph2V. i�'0���;��{&h���1�C�)/��(��~�шPL��o%�R��f�l�)��cB��~e�v�y�/��Zd�z_��xv�к6ha�°�c0���zA!�����b�a	����V�0��s�v\���O���S������{�O��y�<��1�&�`��+A�ϧ�07V��\�M�M�k�>ӻ:�N4 ��k	�s�dfg!QJ��іTb=�a0�L綛����7b�`,��Bh�E)�9�T��Jh���ʠ�"OH k; .`��{� �B�V�C�c���a���9�� >��qi�-A5 ��{Z{X��Cg-fq���KAZ�|��4�	lg���:��l�MGN�"�9q	LEN�����	n�FG�|q�})fX(�a�n�Bs�����vo�S�
��1��/�C\�};��ɟ�.��_�l�,��r޻``�.8�3�Ƭ�9�- �zfz�./r�� БM�g��<�.�X���z��V���U�+#`��Ojd��%�ÃY,]c��C����۸U�`N!��TF� 7��g�H�}�"2"�b?�]gT�w�$��"�zc�h��Z�Њ�9�8�R8�Ҍh�Y?F�n��S��te�$���J9��T��-=kE@�\	�Mփp�d�q\B�2pL*�$;�7�u��͎$s�x��^3'�\
�%��N�*Fi���}��>fR�i�'�}l�$�!�fF`�hH�;���Y����x�;��s����~�-?��8x�<���'=�����N�1S,M�v��w'�����Z E$ L�%^jV���*��V����q20f"�U+(n<�8+'�;��9Y�Ƣ�=t���X�Z�`v�����A��K3 �0,zW\��    IDAT�[g�܁�E�4 �`���sS��1�F�ڭE �x�� G�ƍ���@�0��^&�&�;L��5S�dJ��Eo�����gR��'���${���D�+��5l�B^����D��Fw�����/�0��7�m?�a�}�Ҍ�o|O���qr�
v�8<>���i�v����E��Mh���p�m���J�%���c@0�1ͥ�ixٯ����~S[���T�@Ș9~o�&�����¬���k�R<�ƫ�������+i�VjmM㭵q3+x��a%���7�Fv��_��U��R۾����쥋x�K�é38u۫�<�8.��Q<��Wq�0L+���ڂ{�mT��jև)�k��ֹ�������r��>"r���7�z��%=�4�o����R�PW�G"���d � ɿ�3�B��1�8u�DN��˅���>X�n�h����ג��2��{S��]I4�c��ޝ*d,����k���<a�����w�ܣ��hn@��w��8��_�@��Z�mv�T�����v+x�"����g��M�\����i2�ݱ���)S��kLp	�k��{a��8�5TAۦ��`/��1!�^\P�3v��j�Sp�脬w�V�J��6��X��_ɐ�-����9������S���������o'�c��y?����7a���5��9aI=fMef˕)�������]q^+ckrl���%��~k_x������loHR�]�n�n{�{����e7$L �@+e��Hhl��w��P����`���a�\��M�ĸܵ�Hn�
�l���u�ޟjs��`������0=���g (@׿��8�؛q��P�	���?��O|g�1;3�=c�Z�~U�k�}y-,$Y�T?�D����؄�rj�$�e$:Y�������Z}c�Li�D�����5�M�a�8�nU��& �1�4�!t�8��~����*�����٘00U&d������M��#<e��uo����k8�֢�{t'�8� ���*��{����?:8�ț����G8~��8bB�f=ÚJ��,�7��d�c���S�M�$���yR��p�b,���es����n�ɂ
��?�˺Sq2�a@�M%��m�PG�d���,{9���ar��_]�R��
���}�݄Y�&\�Fc}t�3gn��f���~��ʯb���0�5��<���ٟ�������\Ǭ�Ew��B�4�S����MN��[7e�nv~���T~/�>O�Z���p8^��0n��U$�w���)�SJ��}r�aFo��|6�R
��˘;��Ş Z?J����-���������V#��z�h����H�6J<L;s��
H���)��-��+)S����n��q�� /�s8�v��s'��]�걷�峸x�#�w��3j�k�E�N���{��4xL��<fJ�+�E+�9q2�@�*�%� D���P���~�-.�\9���#s������U�� �HSJ��?�8V5α�3�����#d�8dx�tq� <[3�OI��6�O)e�i�e���{�p��Ǖ�5辇���k8���qj��\�����.��|�b���e۝͡�P��+,��m`���cxO���C�v3��;y�l�����njet,�9�|Q��,�	y�����ف��x�E���Tm�`����\N=Dl�$��������#�S�v��m��6���/uA��br����<�}6��C�A$f���;4��m����x�#��S����v~#��]��X43����V5Y��p�8|�Χ�[��z����2=v{��k�\��Xه��I��"�[� �"�,��ƺG�U��$�vb��2�Rɖ�^�	$�B�[¾��ކ���'vy{�iЬ���.^����so�QtKB��g��?�m���'qj���5:��?���E�Ֆ��$%�<:���'�>��=���lZ�c̽��67kc5ֶ����p�)S�uS����cQ����G�u>@Q�C
�?c`R@l��i<�u[��l.Stff_�O���1�6�N=���|-m�\�mK9�7��������
���|�����~��c�O��������bt~�����<�$T��m���:P{N��ل) �����!�G�M4h��Y8���^_�����N�1)1|�}1Ơ�{�}��V���rK�@�&����R~�֧�w�N���Y{n6����Wq�����'ޅKk���ů~_����`�VK���h�q��Utm3�wS�S�o�P�I���V�*?rQ��3��v�m�ڭ�P�m�٩v�a2S8/��2~��j�k׮��:h�Ѷ-�]�EkW�/����=�~ҽ�f>V��W����8��v��Yc��E&@gPSs�Fg�ʘ�[hww˗�a�q�Ya�4p��y|��?��O}{8����;p��߆�[��+��GX=>>�f|��1E�6=;,'Џ��ks��Kc�:6�6�)�k�R�#�+k��պ_�W��Z&�'��&�h>�G0ȝ��L>z0.�<t�;d��֎)nazv��@5`6ѝ�u����[o�S��Հ�a�
Vu�d����cc{���1h0��3�� �O0�l�oM)S[9 �51�\�.�<�5 �֪��,̦�8��P��c]~�圁F���Ņ`��[p������;ѨX=�i|�w���2��]��5��0S
Kk�&�V7�w��L�]��s��j�'Z���V.N5��H� ����K�=���GC���.�����f��(�4Lۣ_ �0�K�@�@V�j8�����(U�pj��$'�{ƢA�6�U)?o�s��x�\��)w^>|�Y2�&���c$�]l�F��D��0W5k��b��a��g�̜�
�C�ó>��)���KN��u��M� +ԧ��#҈)�`(¦Om첌g���m��;avGR.Ui�T%Nj�Od����y�.sa�X���vк��i��X�`�M �IP�G��z3��&<��M%
 ��� n�5J�5L������������\{ǟ���և��z���pߛ߁���˭�����Vi@
��ԍB�<�W )zM��:�a�5|�q���*���ӎ�Y������aݬ;���8���^1"���^�|�?a� �{��[��{0�Ӟ�4���۸P�g�d��x�Y� hjAp4+ui��[ZD5�#?+�#=�Ky}�Zzx&j,�MKMS�׶eL+=5�G>}o�3ہaƊ�Sg����ᶷ<�G��X���O}�S8|�%���=4�Ma#Vj�H�p�p��0w@��DlQ���"�=F�Xh�A�`5k`n�����vv�X�ccp�8HBd��a�� ǢF�Â��6'��Ɣ�>G9�Ssdb5VJm%;�3����Q�E��j}�pL�m��LYQJ�7��|��8��P�v-��8R+�4���,f��ƬW�zc]^h�D��8?�Z+cV+fF߯��g�M3�L5Pk�}cq��gq��t�����x�ïÎjв��?�s	��=6����r��ޛZ��fF
c,��()
��<
4�h�&��ё��.�WI��z�0��r	�;װ�tҋ@!J5�:Ǒ�kt���{�̑g[������O���2E��fJ��`MVCA��y���pr�4�A8��/��_}��4��E�
L��|�HG�'���K�4�ߑ��sgJ�k��Et�,�WX�3v���.�]�N���Z�naw�a��Y�S^>_��S�tl����q���v�p>�����϶��pB}c�&�pVޯ�1�[t�|(��c{�c���
��qcKW�ʆs܄����sWð�%f�ŬcPg�֦��u�sf��9������-���;Sc�hp��QX�V պ��n�3�<�]<��o��?�����ӛq��Ǳb���{��O���P�G̰�tKY'mu�ܖ0��H�[s&/�Y
��o�ɣ�p�a��e��7D�֤ڜ�p2� �~Mx)}���bR��D��=C�c�х0�p�a1՞���&D�b):5�iS�"`��n���*죍��ZG�w���hp���s���a���quy�ٍ����!���8�hp��.�_ɈʾJg��3#(��y7�3M[��3X�?c�+�����i �`���V��y�A�ػм��xf��j}���N\ٗпm	]9���Y�m%w	������N�-�$e�5M������?F$��-ǱF���M�}F�nml}'M�u؇s1`��eY�k�U�V8k��0;Ѱk ��i� 2t�=�on��q�z�����^��X��I)�3zN�����B��X?�e\����g.`�{;��8辇pa钳80F���ΰou�;Տڼ+۬�1:�[Ei=�I���G��JZ�m�ڟ��G'I9!;"��F��q����c� �*"r�,#y'k���I*�Ob��i��Y���&�����Ci\[�����G~w��p|t��Z������W��Y�r9�O���Ҕ]�p�of�����9-�c�}��2@�C�p��ZX�̱X,p��8�����'���?�?�����B���]�ʌ1�қ}lQ�{�I�ilk�����:CYW��P16���"vSQ��`���g��>��\��,���؄�A �cP_�8�mm����	T���R0�Z��R�,��p�M�1GTG��m���<Å�^��\?} �*�L`7�<W+���T�`�3j`WՂ��+t0��[��,��͗0�g_�f��������Ƶ�Y9I)��@Wc��}�:6���mل�M��X�JY⬸.�Zd�5>[�}Y#7s�H�%���R�c���Ҁ�A�M�|m>=�IK*���f���6Მ�qJ*�� �K��=+\�-f=��}��hϜ���'�Y<���>��Fk�?K�vd}v�|*$S*̗%�&��1��v���Pɹ���г9X���\�z��������]<����a���q��bi-�߀1]��FdƎN�Y`j��o��|�V���&�������T�4�1x��%l����Z��m��1�l��1X��G&_2�C:��C��:�I���g�����]��"�����߀�1֍[O*9q&��9�m��<U�Vx3rCm� ���>E��sl�e߃Icݯ��^��/���z
�f���	<���n�V��z[k�'n�pȡ��!��ܷYOSnYwM`u`(�	�@�h��G�^	�ر����!qVc���z���mN{[��9-^H��<s+Q0�i9t������@2���0��9��L�4�m��8'F.�ݘ&R{ǲ�j�v�9�w{�]x�{�N��(��c��.����}�i̵��34���K�6�S�3p��Y	���M�[�I" ��}cv�`�O3s4�1�Due� K�L1X[k�(FC�'G�݊�o|3^�����x�2������q����nâ#p7N�$�o��IB0F��b$[P��|��l�6�ߢ��h$�荽+�0Ō���&i�n��l3ܯ	��Q֙����P�>q���ȶ%��;X}�^Hw�P ��>��4蒗|���N߆��^���{�?��g��w?�Q�U�kV;U/Z���ao�D:*�i)���1��� ��Ō ��gemqf��������bv������5���`k������ֺ4�j���6	�@�ZZ@7ͽr]QF��30�и�M��D�cD�đه�^ �2�B��bd}�kZQY,��\R���cZO�;g�����o(���_:\%8�zL�ۆXL�m����&$��n�=���,;ƩW��}�O��Q�n<�����7��S�awwL��B�~t,���F8v��@�7�"ʜ����}�0�
�������}th0��~<���ٽ����_ǅ?�]\���p����s��Uu�����,%�j{˵:�:�f9o��i��Z��h䲔��n��D����c8�%a�_Ã�]������1���ڙ������7���~yTUw�c޼�0��   $!�H�HJ��%W\*�{m���7��������ՊK!J")J�D< ���p���xW��􇬪Ϊ��~ �Q�^ב�?3�W���v|}#mч�s��秐9v�����O��я4Ǧ�|@��[ec��=W����%��sB+�<��9�Z�HPSK&S\9��?�K��&�_e40[[㞏<��'�0��&�k��eq�cs۳����ۣ
�pH;7A��p]�8�f��0gDV��غ�9���3g�����<��R�`Zi�R�cp^b��#/s����Ei�� �C)I�i"8�pk�F@�suk-�BR%A���> ?�C9�q��Rz���GP&	�V��n|T�@*IQ�8�1��b���ul�ր����w��u�*��p6dL*���;�in������ck3��k����?�n8��c��O��"�\DS
���0x�ϳ�a�@�>�N΂F✿j�DԪ��;��bl�/�h6cS��H-��H�� !YS�q�l��r._#��������$7�a/�k�.q�/������ ��ز�Θ������L�2���i��h�%�R|��J��<V�s>�����
��\�}~�J�i9��62q��{��%D|~���E��jU�g���0�w��Y��Tkl^`�Gb�R�����Ӿ H>�@� M8N4kY ���CӺ��4"����6`�b�{dݽ7����{~��o�
�P������7�:~-��ߊ<����3�ua��o����cb(�b�l`fSdR"��c�u]=�I������x.�M�]�|�.�VH,����*G�;fɀck�$;��Js���nmc����ˌ/���lB6ؤ��DLQ�@��:9��cq���^kU��eW{������R#���f�J��%%Z�Ֆ~9g�ƒi/�O˒InP(FiB�
�rH�VV�VT3"0NR:0�׺�D�I�Π���Pʏ]*��%�T���U�7� \� ���y�\N���d��qeYѣ���8��w76p[�h��6 ����\i�
�{&3�lG�ֻE]�8�e�K�;�ɲEu�~&d�&I79?3\���q�}w{���}���W�\�iY`�֔� w9*]ܨ]�Uf1�Ug���)�m�������c��2P妤0%NX�����G��ƅ����:��}�3d�mQLv8q�"?��/��?=Fb,i��Sgdݚ��������J�]�����<t�j���l�Eªۋ1%}�1���ol!1��eg�ݠ9������)��1SPG���8�/�5sUe>�B>5��#�����R�"���_��Ў�~]���Ӌ�b2�rb}�������"W�~s��}���g���ڥ1[����!����ּ������g�b���a�.�]�� ��E	ŌK�>�/�fw�N��'�c7ތf[2=�0)3+�:�$��}TDw�q-��CX����{�֚$IPJ5���ºb��hZ+��ss-�q���n���:�P(Ŋ�Xt�N��ڇ܌%�>�w��Q��
1'�aD�X�"��"�p�ɡC�]�z�����p4����^s�{�e���l�����'cp��z�Q�K|Cas葆¶�j�kR��NJ�����#§.�:0�Q�p�D�����)eiq�d7�ŝ��,�]g�1c=?��_~�7��wȷ�"s�<�)]�u%�έ��5��n�g�`�%�ٻ��#2}��p鮿UH���eL�2frU9��bLl����w�+�D���8y���ǐ��p�e��m��Q���5��!�q����:�%�J'u�&Qi�	��e�MgH��'�!���_�s_=�.7��Yn��Os�=��ۻ�@e�lc��dC)�K�����Xqε��%PLl^�0��������5��~��$��nč7��Jr3f�R`�Y�ro���2��L(���~�k��I}6c0]�\eDm�Vi%j��ۧ��K��^v�L׏~7fI�trn,LNщ%�f��J�9�&�M�l�/.$������A��,�ޏ��>�!&���>�#��.kJ���Y��
WA��i�E7(Q    IDAT��E��`��|�=*������~u1e�s�����`E����,˰F1>����G���%/-�f����^��_��{�k�C0���a�S����2/ˤ�.�֝ﾲ
�tϦcA8~��ZW����Ga�����X�1N}Pw�K�����������F>TiyƤ��=���x�޵��a���j3b_K�"~�SK�1�tg�F'&�����x����ܷ���ŗ0b��]��O�噳LP(aH�%���j�I�V��n���o/�a��|��\��k�e!w1Pl�=�S���?�r����?�Q��f&��
�e�Ÿ�����!>֣0�}c��#�Z���k��-��p���B�}���[�v��/�kA���}xSv9�����<�����fU��.�kc0�:Þǆ�"���Ήza�p@��ǒ��&-�2�r�w�b��s8��7�ؼ�n�hD~�m^��7�{�)!94���`���>
�Vʤ�j=���X�K����QK¸S����EʾX�~���m����KO<�+�eŘL��`�u�4[Õ�	ISo=���hL-�kW�Jٱ���'��[~5"�_g�p��v�ӹ���c����K)I�"�
J�d���}L�s0h׏��u�^Ex�r�C����6�1e�#�51��^d�c	��4�%�O(�q�H��l�7���\��/�~�����{胜��O��~�RhL>EP@���
��#��]W���Z|w]���a��ST�b��g~�䙟1�q�����#�G~l����S0Pf������>b_�0�]�_|tW*�ה��p]�i�����{o�v�~7�/Cc������Yi�!!*_��;��c�� �@� @�/��\��w��L�������މ>s���<��G��N2�6�����mg9ؽ���ۼ�أ��z-�BH�NQ�R���ح\ڶs��u��M����~б=0k�HWZ�r~�n� ��\�Y��!����
{�iJ9���ɿ��$o�#$g��ԉO�Q�u�&�t1�d�:\��w�QF�9�2�]����
I�x���G��z����� O��{u���_sl$�y��j�Z�v���\؅6�	|��	J|�,�E��l���9,g9I�aeB�
6ӌ��e^��_��_��F:q�#��=��#��mv���Pޠ�v��$86h�;�n��g����©]�&�i�%���䰴Gq�M~��_a�ҫ�ƻ�4[�>�4S��a��V̎n�	_}�%T��������1u�5Ax�K���Q�Z���Q�Ƙ޹�eY����gw:�t��?B"���(-�@8k��Yth���%�QYB�nPM�PΪ� Һׇ���י��K��6A�q�]��&�ݷ:t���#��]��[et�:�����?%��+�rLj�1Z�%u��eFA�4���6�y�.����u>�����:,�Ɓ�8)p:ũu6�{?���g)��Q���5��w�U0�g
I�h}��̦h	�������^�Rz�e�˸u�q-)����E/��o���(�������>��Wwآ���O�]�lKꥹLr��.#ў��b�Pi�����H5�~tC�.�m~�"�{�9X��S6�C���SJ�ԂV������]^���	Nmmq��əG>�΅�\|�뼲{����{�87~#9o��������������[�B<c)Q��m�UܺD�}�����F���P��g��{���'ٽ|�a6�L^HȂFu��]s1A�~&"gw]A;�_cc�߷���"{A�v���6.hI�`��]�K���G���Q��}o����P�G>QB�d�ĢŽ����9����Y���C>1o��?��EW�����Ω�(Na��X���\����|y�)�:��t�2?��י�}��c#�d�+f�c�C�4(mA;HT�������1�]˂��|Y��7wH��)�R�шL3ҍM������a4�$������|�Y6��� ����p`�TXRm�䇨�n�h�T�%���'6w}@�X�`R�e~�ݲLJ�G��.R�Cr�~��%O��<�����T
�(���&c��u��UG�������k"��.��B�};�[?c��f(6WE	��l$�P��d��1����~��/�淿�*��i����q�ݿ�=��۫�d��"݈��0�}cj���A`l�"Q�T�tʰL�n�aY���Ɨy��믱�;n��~n~���q�t��tns��#ײ�׽_��]o���=Pӕ�خ�o��B4)���ڥ��=�P�����Nw�V�u�g��x���q��4A8��^R���4~�~d @)�u%EYVzuϵk>��3��WgC�:��,q��6��h�b(�_��|p��|�3�D
�D)��c����wmR3�9����5u��#�#�G�C�K��Sw΁sHY�9�:����kK�p5E���^'��H�Ag��N���M����7J�V���.~�k�H�L�K	��-6JS�r	���[�)��4c�����yP���[j?o���b_z.S �rƦZC̼�'I3�88~#�������~���3�}����?p�;�`�)JkF�8�p��K	R�S(�|�p��>�n6��4?�
�B����/g���輚��7���;"���UˊG����沂�oO)��U�n�ж�;�.B��R��a�"�n����a b�k�y����f��:-��>�U0�FU3M��k�\��B�:��ffi���R(����E?3Ε(�TuՌ���՞w�,����}��� �}�����!���-�
���˜�$V֠t
B�� ?���s�sz�8�c���3���7�z�+W_�MP2�5]�.,F�
���h�]�_)�ǈL�^'��z~O��HQY�;�0!��D��y~	7p�=�o��G�{�g؝���\ A��	R�"J�����c%o��z��>V@�@V��1#9�</�J�h����]%*�D�ERX���$��T:TR9�3��)� ��AiE����PR⬣^��b�K�qe�tl8��s�}����3�yf���Dcj�.�b�J�GQw*�]��,��ew�J�7���x²Lrx�w��	����ƚ7X����";u=�=�QFǶXw��W^����I^RLf�~��ҧ����zgq��j�>�׊W�e��R+�xק>������������K˫�~��L3&����������m�o�}�j-�m�Xݱu~����UgU�L��b�����$��{}Y�����7�y�UK[���Gc�\O��>c��e��X���-S�H4NIr,S[2�%3g�E�	M�ŕ[�TQ��̷�N��y��r���y��|�������d(�!K(J�$����N^��okB��iA�{�q����"�'n:˻��Ӕ�$Zz"���Qt���qSC��O�����}�5�Ƥ����-O��.��R�᷍�T�X�iX�HW�ѕHb�
U��D�����G0��Qu�Y6���%6a���b�h��kC����"�`=r�K6o7��?��h2��Op��/0b�D��o/�����j\�P��Xh�4�(�P��?z�t9��g���'��qQ'l���ͯr��_c���p���,�J;���ֵmHm%(|�'D��i��-a��k�hua[C�B����SX/CN�>�%v4�G���>&��/�{}�M}�o��/�v��V�����G;�K���ѵ��,�5���h�Ȁ��O�Y�3-s
g!�dk#��!.Q���<}�S0Њ4MX��g~�Ͼ�e�d�])8v�{���O2=vWfcReq��"I2�$k�v���(%��b��P�g��\�\��12}�u^|��ߺ@>�b�އpۧ��R�|�8-qJ�|����D ����F+�m�{���4Q��~u.�>w������� ��XHS�׉�F]`?�c+^_[�K���߬����e�/��_6����l�s�:��_BiZ�c,w܍=uƕ��q���eK0!5���h���Iv��|0��<Ӈ���(�`���hj�W'�N�ɯ}쳤�[)�/��׾Fv�
gNlS3�Y�v
��o�P�J��o����s�N��.���=T�w�X{G)˘�p\1D^}�a�=J��b����ۿ������}�s^-�	J@T��b����� ;�h�hߐ��N���^�e�iJ�e���s��IN]w-��۬��W�Xj�a�=RR�֞�f�"'�d͍����O���8�7>���f_I������I��YtN`�+��b����i���~<���ZQ��
�ٔu7e��S����۬�v/�~�#�WR�VB��
��,KR�E�[V�k�Z���(3��]a �^�:H�c������Uk��C�E�矶l��/�P���.��Z�I��5xc�:����JZ�z��ZW-�ظ�ԭ+K4ɚFZ:d�xkz���[8~�]�)�����e���8�%��Ô�([h�W-��rf�.VЊJ����`,ؽ�6��o�G�ﺓd6ac�<�����ҵ�3%��� �X��iB"����q��(g��s�#j}L`~-D�b��8���n��e�iU�.V�C/2b�����w��[����{��������h,k����6/1���p�xw���._e��զ��P�RR���"�A6Ɨy�O���K��lIy�iN}�a�[�`�2L�4# Ԣd��{1��2c��(!�RڍNX1gu	�:�(������*��1�Wv�k[������'���a,(��0�%��UWw�s��%BO�ӎ��)��5�-���b��c떣����Њ��݌+[�cb�#t]@uTx��|Ѳ�:j,#'y4$�W�qC�>���(g�gS��1[�M��\�2���'����0� Ǘy�'?`��0eN�$;����,��5��kW��Veՙ�U\����+/3�a6d��i�~�X���9�@M���7��ۏ���Ô\Y�EI�S�Y�y)�_����ţ�>�rTF%V_���>�a�G9C�c4����w���O��؞<j���UD~Y�Gm�'��m���H�a�g�T!� ���/���K���%���}�/JK1�p��Gy8%q�v��к*���$IH�`�ed��W~��_�ϘW��̧l�s77}�w1�o�ⴄT�LI6�a�ø.�m��I�k,R��<ᓴ8�p�@� �JZd�����W~�*w�SgX��יe	c[P����U�������.����=˄��
5Ρ6��nn�)��Q��C�o��9@���,b�*�e�,ƹw%����hw���� 	����"���4`��Q9dߠn����ۘ����+?�����LSN�'HC�XqX���q3����뫳�7P��n
W������?�N�b��O~ȋ�e��)��!�B1t�I1�p����f���w���/Mw��+��6v�}W��z��-[[u�bAy�{}.}�������Ǹ�b����UOHJ�4��vl�e�o�l���%��GMJ�.+B�J�؛�2J��YB,&+1�0>�!m�.%�9d��O}�+��;�7^cm�7~�c���OR�>î�1�3��בh���>�C�ƺeq���q��V!D`�V�P� F1+r��e��P����1Ǯ����]�u'�j�Q�+�t%FXd�)\�r�W1�}�:�a���m;F'c4q^G�b���K�k���S�8\3���0�!b�(�9J���󩥫vv���.����"q� �e�#V�""X�1�6�3������v�F�d����ʏ~��X�l6#/K2����'��[�-�ɯ��{�������i>��g}m��"��s?�[_�÷vH�d�Oj,n� �9�ZJ�rR=�H*\��q���g ����1H}�����pGa ���{o�CRݾ��lN��_�,�;�>��E��!jW�91�_�5m5A���Ǿ�,���1����,yYbq�/˒b:[o����4��l�&C��;��Nx�k_�ҏ~�����u�������h���cT�Nְ��"�o]֍ߣd�dV�(3^~������02ct��=I�hH5z�bl�<%�i��*��c�s�kq�ދgm]�\��o�7�=�j=�%4oK�̝A�;���J�LR�&"��?y�����
�X�u��Yb��o>AUhSW"�Z�dK�\+�m�9��:^q�a]��3��8�����φ�$8]�kZ@�M����^��/��xNUJ�
��J��L2�6�c������S���O��}#E��O����8J85"#�%S5��s�
>�L�0T��'B���~��ih۪���X�y�P+���)�vks����g�?un��Ǚ����e���r��_Ƽ�c��5f6�(Hȇ#
%PӒ�K02�
�D���R����
�>a~�znJ�(�ø&�_;���"/)��hmp!�i}ݢJ-�81"Α�»�:��R �5�����ZE���:�zra4��-q�� ���ۅM;��i��ZW]���k"�<sE��(hjKv�֖#�\�3e�V$
%����ÖB� �y�ẟB�&D4֡�D	�
�����Jb̐��:/w�"~RP&����1��xm�8%)
�R�}�0(�I� ���]^�����(�j�;u3����8y�)r��,�Zc��P�b�43R�pI��!�T�/Q{7�qt��I����u9Uw�Jp%W��(P*����)��~B~��t�N�x��?�>v������шLM��{(��Wmx�PX'�&�*^i+e��8�ο�D���$�~=9c��c����
��M�^X���T4)MS�N++{D1�3+�Za� ��q����-�:�1��)��g�
\uD�u��CRc�&+;B�H��@H�LpȆ�V�g5���}�~�/�23D^!Ҍ-��T���wҏ.A�qY�ι�𪑊���]?ƻx�ts����+<��G���`]I^�X����I`W#��ˬ�'|֧f���9q-�o|�-0yHT�!]AjK
�y��������k� �� ��w���͡"W;+aݍSw��ϲ�lnc��t���2�7և���>Lt�^��>_6�>ɬ�yw�����߆0���Q�U�m�!<C��kbg{5zWZg;*��ﺟ�~��t]�)��s��[Z�����~�}?Z�[T'+j<��⋜{��%;s�k�� Ɉ��l��QN�h���4R%U�UIc��я��<-+��=�h�p�����Oq��և�l�|�n��%��a�K�67PI�Gl�X�5�%��v/��S�]�c��{�F� ��-Bo��6�+���m�Ѵ_yw4}��{ˁ k4�r��|�Ӊ8�X� b��P:�\��GD��2?ː�nX��"���ބ�̻��cg�}�5W0{�u�=�J��
�A&zAz\F��������Z|�!�b�p��z|��@��)f����l�� ��1��,���?����W��r��t��)��|�B�F��6va>�TV�~ƬV�"4�������2F��}k���]�b��n���e�\V_wE�ASg�l��ph���>:��;��:�$u� �/!��3o[�*M\2W'���x��p�X�?����K�دj���h=���[�,�\A��K�7�G�p�[��a���A����,E㼶C$��bj�g��iY=�~��N\3T�2��j�JXO���o?�c�I�x�N�u?l�c�2В�8
�N���ZSq���e��9�x����j�����j��y��>氻�����.dtk[�����m�AF1⣪P�M��uK��"d�A�	~TFo좵n]ˁ��k��q�!c!D�}Ͽ�/��
s809�)'�}���n��9b�m^��o3�g��ګ�T���qG�.�˯���u�`���o��NgH�o���o�>�{od_�Y7{�������c+�&��q�B�F�Ssʦ�H��O�}H�(sK��q.z���K%����v<�W-�Jҭ��Wߺ=ʺ�ǵ��c��YGU����+k�(#aE;��dRk�����_g|��.Bj���p|}�Bx�Bߌ���&,����O���
�Q�:��\Qr����){    IDAT{��O��[����>:�Y!����:E�e$I7r^�h�o^[0ZFLd��/$�Ɓ-J��#$��b�p���~���[��s�Ïp���0��$d���n����>�+��G?�D�1�1v�~}�����儂o��B05��	W�N^� �׳]���o� nގl}��ѬS��d�ٺD�s-U��ۇD��¿���71IK�pF�U!�����҆�?����x�@(�3puoLv�����=��\y�����b]*DQ2�'͂�t�����^lA7�;`����X����`���}�r���p��m]������3O��5�OI���k9�s����q�p޺a�[�>b�m�<Bi)y*V�s�{	�Wؗ:�DW���X��@|/Ş����c��-L�����J���#��R���\6q�=R��vT�FU_�1�������8���cs���W�z=8�Ota�Gb�L�����:���T$l�}?���g\c'у!Z{��ٴ�̋H��ġO�m�E��f�b/X'��$6/9�
���'���w��u��w���x'c ��`����*5o�u��1t�����'�@%�$IP�F%�ٷ���Q������I����?�:j�Ҋ�y~��j��>[�0�]��b�[5ϟC-�F�Ჾ��s��׫-�z!��)��a��Ai�㡇��� �f��r��3��dJV	]<�po����18���ژ(v�����z�Z&>Fw>f4Xcw�0�o����<k�O�ؔ�[Wy��
��O��X{@�Ǡ�ޥ�x	���>�H_8پ4�}p��c��K��c.5�ڭ�u�<�1��I	ZK���*.�/c� (@׿b�����}��^���(���&J�Gׅ�;'�Z��������Z��ma��\���얭���+�x��^�3�����;)G]�B�f�Ϊ�S7m�s���x�k_%y���\��������%#qY�N�,HӔ�t�� ��FG-�p签G�s"Ek� 'Ha9x�%~��oQ��2�����\j�R]�	Ga�$J�=�W���H�.���.�އg�m�*���&��Llm��G0�~r��R������̮�6\�xc��(�}����0�A���g�iY�:c�V�A�e�lU	��1�Q�7*�c��M�(�b��k�0+8���y���F�J��!u�B!�C9|jZ׿��~�NB&��[0��]_--Ed�&r�K%VY�KJ5"{�]��8˄)�._ᵯ��|�K.%�K֫��;� ֐�粛j�w>z�[��\9K�{�t�񻘼���[�>�ƨM��!��932D�~,Cl�;1�9l�
��E;�|�fW*	$���@eY׿Jҩ�XK�����5%|�t�:��j���[����үVB�%��m���p�e��7�������9ԴĦ[l��>��7�oJ�+�	���yG��;��*F�s���}$e!��8rla1dL�cc�W����*6n��cﺟ"I�N�NN���d���^��-���w���t�d6��yN���>�7�7�i���e}|�����:c�g.�����p�Ǌl����Nc�s�&�Z_�1G��vaNBB�7uQ�"�@Y޷�5���� ���Di=�r~B�C:\�&�ǚT��쳌/������`V���}��Dy��nT���;݃ZR{E��p������#-õaל9��{��0M����O~��e;��S�-4ÙF�3�,Y��A�Q��q���QhL��[s�\�6����i�b��49y1m�sm[V�����/�s�ϰ�i���\�c���FU_�~oJn5�`�	�3�n��QJ�(�2�/+��mǐ}�r��(�.E��q>��u'P�x�;�BN�l��[o���j��Y�����1��t��g���>�5���_e�-�t�!�����Ll�e��^x�\:�Y2$��6O�����:]ۅ�cvC�PK���fa1A��`O����n�����.�ע�_����Hp�!Rz��_h���5��Y���,�x�� M\i�JW�y�&�������:� Q>#]"e�����ʨG��
'S�P$�D��I}�7�Rz�d��YI�[�SHBX�H4����8Z�j�[5L�!C �%0+n�#��Pb���O}�;��/~�X�2����K!���Y-�HKQ�؊�QJ5y�-ՙ�h����s��?�w�X��0��#%%��h���`M%I�� �d&n`@����in��r�G~��xFy�e����}�*��l�1��k�����IL"��2,%�̘�uGǹ���]�s67���['F@`��|�+���-�\��ȇ@���ZI2��Ɓ,)UN�*I�`�g)ؗn�2:�)5ߚB�P $��
�"����� �[>���&v1�c�zU��P_�J�����v���T���_����~�xfT���{�2Od��Ü��=)�A�� D�'8t���U�m�Ъ�܄ ����#5�e�Z�x Zq8���i���UF�5��D�H�P��7��ؼ�F���9OJ��cY��>;{o#F뜾��R��ϾHve%'h�c�U&8Q6���FV�H �~�i+<.T͜{,�6.ʲl�H=߿ �M+��D
� �($8�/\Aek��vN�r���+\y�E6�����pS�3�
�ʗ�v���\�N��x�s>r�Td�(�ȴO)���MBxC��	
k1���
g+&����j]y�Y`-��.a6��@���
��TX'�U��AYz��Tg�i��G_�l^��2XJJ��w��_��_�$�H�3�he,�U�<���Y/��߾�m#�Ru�k�����8ι&p¯Z��A�>HS�0�HuJ���?�������I�򐗞x���|?J�~(��6}�`�cR�a*������R� ��!zu�`0�=)�=�:\g��;)8���s��{��t�K�z�7�~=�1���p�C�Vm֒��l^ �d����������y���.m���d0����9�5��О�^}�@:�� �sf��(AST���&w�Ʊ9)�bʚ�O�(����x�H<�#����r�j�׾�O�+F�0\V�~(�����[g���o��gm�ߤ�//����/{��%/wq��l�q��Sg)�c�ю.9��1	,��kWb�>����|+=�*T�lZ0�)�x�������N^˽���\>v�K�h�I$�,!����]+���R�Y�;Kg���d3�����k6��/?�-Ƥ�6ظ�y�q�`�fqW�欶1��c�����I)��Ř3#Z��� §.�zo(#_��Z���x�M$��G������sM<��B1Dۇ|k�S�Ď���%�ֻ]׆n���[�U/��e����"(ϵi�m�3K�+ԝ��q�m�l����=�{�
*QP�diU�k��h/:���0A�AQ�
�ߨ�eG [-:��7ƠF[�\{߃��7s�N��>�Sfo\d�X�1%2�H�18�Ш4C8�(}�3kK��f�a��㜼�Z\�B��
�Ӂ����9�I�1X�ΒI&}4?�-�2gZ��Q#��Ր�g���`@�#�$�T�n!"�!�&0N����B8�fm�H�-f9B(�
���y�3�����:��%[��yD;7�T�[^�݈
S����m���!
�1� \������U8�rq���x�5�ay's�m'��:�l	02��0����������(�7ݍ��v`@�[�8G�q#�ݨ���[��G�v�m�:j��&�/��!��e����°u�v���>�0Ô�D؊xҩU%W����u!��^�ٳZ{�5ֵ����1¾j-Ş�̖��Fbm]�>hXH(:���I�]$�E��M��(�Ќu��pP�>!Z��H�V��*�Tir�+q�:~�s�N^ì8 ��:���&��Dc�k�8`1�Á.n��nY (�6��:�� �t����O��ri�y7�a�N����=�c��)Z����,�� ���ɤa�2�8���a�����/����Ғe��j
c�N���!k��J�	��	�1�)2��h��՜�c=�9s;o���1�0t]G��6~��p������7�}AlO�1���_|w~�v͙q���܂([[,������a�I!�<`Om����^����Q#�YK7I�	֕��C����e�*Dj[��Ʋv�inb��.��_
A1˱�J(
C&Ǚ�������`}�4w���q͍8[ɀ$��Q:j��/���}.��v1LP�*���ť���'��Oؾ�Nnx�['+����hvA��"��K���B��6���F��վXO�.؏z�c�F��R���d��;�6���XuY����:�p�F6�L������lG���}/6�>��(%6Q~�k�E�p���F���r涻�"av�^��oa/��@	��ҕ/�����N��tԈͷ�m�U��6A@̳ӅC:XO�xKIn�ݏq��0�˨�_���s�b1P�LL����)���k�JC*Zz{����,�u�ƕ��?��x�'�����S�M$i�V���s�t��^=-)*D`�E��5��1�D�5.�y�]�������[?�G��n@��4�-��~/���"��8�6tL*oI.ϕ��v�/��[���5�/:?C�L{;�ƜHt�*���^��oR�)�fG���u=�o���1�ʰ6,[MkX���ɣ�X��
2���:�<�0�6�^|�G��O0�<���}����:�(�8!	��hL+|��#��]6G��P:o,<�a._������d��'��� �F���&�R�&��QK���[w�C��o��E���~��a�?a=^>���3|V�����Mb���$��u�{$���S��O:��3=�Ѷ��~�0�w�}��~� ׊���*�dB){�fo� ��^~�7��8�����Jʬ�s-f�=NɾA(nޏ:f���\� F�"���z��J�k@|ԥ�SCv�Y�[n�(^}���럒��I
���'y(�a�T#L���py��
7Lɇ�r���ڒ�Z�`0`��&��$IН���$ܷțw\�HVkJ�	"�0��Ӓ��g�����?ñnc��Q#Դ�,��1 F}g��{1B�l��U�X�Qd�Lb�RH)�^���v�W;�z#t�����l��B=�8�Dx�>�����n�C�������M��Ǹ<J��� h-�p^F�cc�>�.�cߖ�!KR�p�2�DHP�P��,����o3�<��� ���2�qŴ�4EÉ��k��&r����0�t!��8#k��@�u��p�=���M&�M_��k�'�65�_U�i͖�C���B��s�����L�,�V�,����E�%z+�j�p�IىZ�<w�2��}&�0�q,PI�[rC��Pme����k�3�i#����)q�w����0�a��9}��$kC�@#��L�k)�\^��p�6�9�	�6��\�h� ��I:P9����[�	�! R�q�����?���&�����_断m�e�]b�(�t$��R
�4�L#�CY�2%�Ʉ��Qf�r��6�(L�)J��C�xJf���:#��UsT_�xk�B�VdIʬ4\r%�k����!�>�!��M��&��/��ޢ�'d�-ݺ�Zf߽[�}�@���W�~,�>�ʼϕ:�U���l����j^���a̍���v�Q�Z�eG�j�k�O��i�3�8v�Z��y7[�<�����������D��(�j���*��V���y ��49J�<J)��
�F�Ή���w��q�����G���OP&���Y�F�\�1uε�U���#��X�zd�(.H�V0q�M-ї��G_�o��*ɱ-N�ykk��l�a8	8J��>�4ܣ1�4���l�Le�^��ص�.Zm,�}}0�[Kι�V#�>�M����plmKʣ�{�aX�N�~�}yۥ�۟#��H�9/i��Q���e��ׁ�����N�9��~�ַ׹Z�q�ܫ��0�%��C�u��5��ķrD�)j"_]�}7G��E��}`ij�8�tM��\��?���1�~q����]ʽ=�����)�$G^U�aV�(qX-qΒXHg=-IJ��7�͸R�ɕc}}��a)�T�([cj��=����P�cR����i�c�ָ�������<r����e�?�(/��"�t��O�sy���&��n���M�}XVտl_t�z�{b�t�R����{n4�F�a��Dk ;}�D���VB�:{�66ή��������շa�"��u��<�Yn��@$ل?��,�V�Y\�a�+����R"��ڐ�tڤB.&6���U
�.q���^�H9�n���?���k��Kǣ��cЉN���օ�gmsU�?��
��1�4�����Ϣm�ю�kOq�����mE���"������a�{
b@����L}LqۀU�'V�o�������3�Ԕ�^��pT��Jzeτ5�����,@Z�V�4Ѥ���g]��(�\J�R!�$Q�4�h%�?��o,�@�3�Ki���y�T�|�Rp,^Vw>�L�FS�P��9��Q�z�����rM��I	�Ddar�L��2e���8��g��?�G^����QLC�18<��*�k�Xg�*Glip�A=��� W��~&���|G�>�~�5��mU��J2kPVb� �!��m�������k�7\�� #�<�7��%R�����C+��^x)ӯ?g�$NH���4��$R�TIo�"�J����ۂ_o����7��Q�7���GV�L�#����C��8�&��0����rm���>������#��1J�9�9$K�W��y����]a�x�u
��jMV7�����}��.��+p�JW%*�^E�'ՑH�&s�}S�����a\M���N:��|�^�Q����y�<����F�O�h�%3��rU?]�����bh{��.a�LB��8�}���N�]Cy�5�N���s��7ٻp��DpX�KHtJa�v$y%�����C
8����sp���l��6G+M�c�8D*1Xd"�U����>~ɉ�Ҕ�ŷ8����d8.�hfJ��$q��t�G_ð�7k��	�%�5 ��V2{�Ϻ��O�h�m[!��	�l9�3g��Lr�q�␗�{	5�c8����La�,Qr�u�C49<��Т}�$��rRT�����|筭p�B��k�1`��:oI�*�����<�sBa̰Ls����$J�)H���@��ǱBb�$ϽP�脡6�dW�H@`EmF&��W8~��8���H�
Y/�:V|}&�À�]j��BW��'2\<�����ͤ�uYK�ͺ�P�P߯�5t��
�kC��Ln+���ӘB0��k��s�2�J�F8�(�3�m�G$�`5"��޽�u�*�RM!(�p8�ɔ��c6o����{/Ce�;��Ȋ)kـ�����F�����{>Mr��~�:�̛6c� X,�0 ̔� 1I�W�,�ږ,W��*���U�k\e_�%�JWW�E�9�$$&���X �����8�3�=���ꚙ���sΓ���,!��|V����xX�17ZC�f$h�]����y���h�E�&\���ÿ���.qh0)����;^��8}����p��ni�z}ĥ���~=�Ei�g�T;?�h�$j�EMw����x���}�5��$^r4�y�������E��$3ǽ>�����G�ť"cs���o�p$3�ҘV��ks��؆�A�o��yۥAo~g�Q�p��s��������0����qD�6B�`�n��p�4�ծw�������.�@>�qy�61��|��Ͻ�3�c��
��C�W���i|�`؅_�㬌P˻�-��*w�`+ ��-��.]kՕ^o]t����rDV����e=)�p���\����uD]?��s�] -5�T���cz;��u�a7���K}�7b�t�z�q�����G��͇�g��L��������f()^��T��Nz�$�N+�2N}��~U?��6�!��RQh0>CyO.b���{sx�Ȍ��o��w�� Q��sh�NU�ڭKa��}Ȳ�Y���5n)��rG�L    IDAT��k����#��|��gd������?���;�2�&�i��:B�}}V�.��ƻ��]Wi ��Yiqt��Y�I��?�+]����y�ꈹ"���U�}d6]��43֜�Dq�g�㕿����*f�}��ğ���ػS0�:ĝ���ڢ�v�xm��&�]��#:����C�EG��N�Eu���+/p��+�������|�;�3��-R�9�<�(|w��.F�=��s5��o�w�c����`���1�LIU���76�z���(�џ�E/�������}8���S��ӷS���	�3}���=�}�+��q���N7�l�-:7�.�����B,�*��z��Uȴ�і/�@u"���ۮ��Ϯ��H�(�B*�)�?�1�>�$~���";��b-��N0��P"��w16]�w��.�T�t��S1e=��̊"�v��Z2����3�|�in{�� ��?�\��fc
�R1��z7i_�]D�!�ղ��.�4�Bc�M�cɭ�;8�=�������Y�pw�������92���$��D�M�n��_���&��񮜣Vݫ����A*�$�:�܅<���5~K������Zo�}jê����}N��X�o<�u�����)�N�$�������䥿���Pn��ξ�������ܙ��#v��x$��O��څԻ�߭�^Z��ʰF�'���͗x�;�b��3�����F9�Nn�K�Pޕ��.�	Ⴙ�����ص��qU�8�*J'���FJrDC:���2������~}��"�0Sdxo�:B��\'}�l{=-i_D���T��t���i������Z[QӘ���ƷMc�EY��{ėO��'a.I��^;Z�tmξ���=�N�M*K��~��j[�w�c�ҵ ��/�����J�'O1A �/}�kܼ�*��$�8�QJ��w\uF�}�#�sdQ��BN�Y\�ǥ^ �f�kN=�>�>�0�.]��+����A b|��q�+���Aγ����V��W|i�������S���5����������8���Q�1)S��-.~��g{�tƥl�d}�a:`:���f8���J;n�o�K��*n~U�]����\Roe<Ww���Z�ܥv�н\,���%����\�����u9W�!�G�>1��`�M��ï��W����X���o��<��y�X�9K���n�uW���`�oU��{�<FF��L�у�X:��6��l�J%��ĳ���3��zH��.+PN��P�+�#��}ޯ��QD���t��?�>�/��։S����9A�4q����9�&����{]�s���y��:�՞�/1�=BO=�TH� JxWa�����B��β��j�A,��T���~���X;�[;�K[J�k�7�8��R��Ou����A�q�/�{1��)��!��	�X���9��"�x�VP�t�s��>�E��/�*�Q��}�ԯ�E�x8������k��C�%kv�K�����G�N�|��8�lc�x�����WI4���N	/���Ň��3���?�Y>�V����y���=��U6"M�,F+�P��DG8�\']�B��mb~U��k�=�.X����	swۖ�}��~LE�_��A`�jn�B�+m���l�h�K*i��.�A�:Y��3��[2)H�60�pl�=.|��y�k_d�w��>�q���?`W���#ȝ������c7\Vk�c�?�|�BƹŸ�Y1cc���K\y��$Y�>� ��z�u���|.���=��^�Ҵ��o�}k��=�Q�#�*$j��\���~���;2ƭ���i�B�V]'�]����W=�&�� �}�R_�s�;��1�=��F3kC�*撆Fl�@s�R}�vS�/���GX�L��)�C/��mB0�.��A[�m��P�{P���$��"�B��+�t�G>�I��{�5$�wP�֣�[���=EQ� ;R�$bmx�2R��zoI�Th(	Q�:NV��l;ǉ'�&9~��t���mn��Qx�(l�p���s�A�*�>g>:�AW��U���!�s�+3������C�Û�;o!��9����H��9�Z�3�M�r4���,�� ui�*<sՇv���w囯�S_��3�>����/����]k� �G]�/�M5%��~5K঒x���O��q[Қ>��k���y�r�h=���Qٔ��S�H㔣^r�K�;o}�ˬog䳘���y���g�s&�M�n%������X�1Z�}�u�4��T�o
M�ϐ�`0�ܼ���<Gv�mf<p���QD1F�Jcr�^���Uvk���������������0�4ki�o3~�u�w��9��#�t�ۻ{�\)��J�� �}��E�&!=R��	��b.���&�u�שg)'KW�����N�8��k�Bi�b��b]��M���T�V�r�w�`[a�\G����:�9�(��4����v��^�2<@1���ܒ;���~7�CG�	o����n��C��8CԎ?�6��/�>[�6C�W��h-��~!,��!5S��C��ȻZ�w�WL/_B[�d:EG ��H��&�6�*�G�ۈ�B�sX� ��|7�~���~ ifܾ�?���q�����h�I"���pk�@�llbo6	�W��ޏ�3��j���>]k�`����B��>տ���;A|�޾�����_ ���u�3�X���t�؞�>��*�2��qx=bS�]��dNa3��>��/����}�u�tp�3��)�o��]�p�d���_Ő�����Ƴ��F+�$j@�w����#���x�u�\�ч���O"FC��H�@X��s���,v�0�1�<h�[�v�1�1�8
뉕$q9��ב�)�C'x艧9|�	�(���k-Y�u҅.����>�l���4�v>�4�z�>�}��ų`Wk���u�5�q�+���c���J��yxU)q���Jy�0H�ё�ySJ�TP�|���-��3]�JR*��Ò�WX#:,�<sx'����,�2�$�,U�:�s�Hk<
�R�K"C���y��(�����l;8���X+֑�m�YC���ۼ�Wϱ~�#3.
T�6C��B#�4���f�$g�<Ғ*���vx�'[�d�$��#0�W��U��@ZO�I�d=̹Q���G�M
n�^�?�0�p{l9��%���� '�0�p�������=M"��7?�lD�s�� �9�
�cl��i�U�
6�:v6fmk�̆,c���qyg��>�;�|ϯq��;w��ů��s����Ø� ����8�8rL݄b��@i��6�Q��aL��c��'2�s�V	9�j�*Cj�p5�NR�B8s���S���1 lM�����sU�^���Aj@*v~y�
�x'�����(�0GB�P��SՑ��]%f�n��1!���ㆺ:��.��L�aWZ
�$$Zᐠҥ�yջ�3le�݉�;����W�y��`M�����c�I�}��gx�3���\���1���
��Ѕ$E��EЖf�� )u�uZ�_�o��'x�/Q�/�$Կ����g]l2%�!ټ3��?�#���2���#d[���txaq�a2�L����\T]M�*
%D0.��-8�T�R��%�0�j_, �@�;r�y�ȥX�ȱQ�_�ʕ/��G���p��1�CED�+��UX��Ϗ �G���`�Jz��Ę���Ԩ(F�/Tm��(�Z�h��Z_��ˆ�Z�*/=s�L�W����4����\P��Wx!dLn����һ��4
'6/prQd�P&a}�ڮ	��FV����s�M�gئOu:/�!R����3��Θ�'�I����g����i�Ǳ�T��>!�e���� �(fn��ko��.r���RY��U����-`S�M���ns��M�R���a6���o�6��F�+�߼I"Q��ޡu@X!����څ�R8u���ީ`���� EG�D����q$�hĥ��H��)����z����b����&��_������:f6��XX���Pe�k�U�	��[�o�C�"E�+�|�SɆ?�+����%��k�9��i�{�qN[ဦ��AJ�
��?!q< B3�	JHf�c-qc�"�<�d�����qq�����o���{�
f�s���|���^?��	b�Ix��'�&����Վ�؇G�Ҏy��ti��m*�=�sO�t|���o3���Ɯ8}�G>�Q�Gh�Ɉ�硎���l\ީ�zW��9��y�t��a��c)&�\�p�;�E1w�}��:��	^(�wh���_�#�׌n��|w}ֿ���*������}<D��z�]���-�/�S��K���O5�<��9�FDX.:��� W��@�IM�V4b8\��%�L�P���'�g�}�o��ǣm��w�O~�$G��3
?f�y|�	@�sYJ�=V��K�z�U�>+�^'�sX�'��*k�	�[Q,X�Cr3������~������~�;�n�$��$sy����;����{\+���1(�E:GQL�l*͚���
d��M2�E��� {�i���?$~�֏�_��W�.��ȕ�e�D���^��c% <�/Κ��(�(��'J=��3J
8펠8%��o�էz<�Y���ڰ��_��"��gҸoH����F�u��rCB�6�HH�d��-�l� ���9����'��9I����_���:������G�i%��DD�Sx�U�$Ju��}c���jF�o���W�"'
�#���E����L�����=���12#�J�ľ�Xu�r�}��E/�2oAE�˧�[��q�A(]2�Ǡ~�õ_���+o�76y����D
E4�Ȣ�n��u8����e/������.m���ޞ��-����E�j�� h��M��\vqp�I�`]>�]�W���"�ϭV�Xn2��DQL!7�)�lN���̚V�r��>n��e8�g9��Q�{�Y�0Eۜ��u�l_����Q[oOvK����֥ͫ�K���(<c2��l�v�YƣSYp��˼��/�E���z�qvn�eGv���k��{%��8�7HJ��($N
���7�kM,5:"������k�?��
���\���9��`�5���
N�����PSȹE����,��d9�M�-�sC���N���gV�߷�b�7b̋�-��b�b�?Ț�gv��}}��8��ɼǥ��[��|�]���6r��m�"!��M��^�֗�\���N���g~�ܰ+$I�1:N�S��_��^Я�	]Lq�و7b����c4��c.�����u��?�0��xB[kzqS#g��k	�9�s���
s[�w�Ϗ-ǣ8�4�͘���^�9�sO�F��
AX���¯��9���Э]���]_�^�(��ei��\W�{�{�pE/�@�쪤ޱ6�Z�/pM)���R���̥tK5U{y�*o�[���ar���q��8�P��enL��M2�<�����{k�d�����|�W��u�"�D�w'~P����/�`�VQ��Lb�n�38y�G�}c���_�s�A��E�-��aE)ͫEң���i_���o#�P��KA�cf�ಅ�v��&��0��x��\��:ͣ��)l]������׾�-օ�Xc��YE$�Ndۄ����39
�C2L��6���w=�1����Vf�5�c0�v��O��g�������ĥ��*m��n5߶��s����{��&�_hۺ�V���-NinIū�)�2C����y,��%���S{���"S���=6Ә����?����f̉g?ƃ��<���!Ɋ��X�3�����K]��۰h�����/$�L h�Y��W_x�������3ϐmn���XK-:�2�n-ý�wԒ�����H(��
M8�F8"ܹ�����2v�,�E�I��$	kæ�}��Y�uN���"wC�wJ�����㫹�� g��e���%��PXrw�0�v���en����s��;	�� t-�: ��&��x�r�cq�ޓ =�:nn��E�<��>\Xb�o,��p��𱐺#\�Ջ���o[p�3�J�9�z��Et�V��'k�	�42�o�y�iT�Ɉq!X{�'�x�X8��L_;O*Z*��b�@����2[X:�'07����s���<#G��>N|�c��CL�A�-4I��L��;t��~�7)┑5�7^ᕯ~uk�42��IӔ|�#:�=�}�}�?c���(��ܼ�����ǿ������'��'��,6׌����>���an�i���q�}ﵟuU�'�J<x��v}��o�j�GQ &�(���������#\6�>�����W��>��S�!���a�)������������%�\̽����c'�t�.]3��;a�n�ݯ&�˼�U�}3��Ɣ9�Lf9J�"�+��{Ư���`��G���{co�G͊|���������f�r5���r]m,��)�!�	�8�!.�&����(���#gY��n
,��m���.��♮��_K�ڂjV�c�c&��N�l����Q��!Ƴ���g�m�w���i�"nr.�3Y�Sz'����\a�eh%�d�_�������&X�JR����N���măH>��	�L��f��0���"�q��`P{V-�D�s+ll�T;3���(�{?w�~G��LY���x�����a�v�K?~�k?�jf1��
��۠�����'�TW[e�"-1Z�B�s�g?��_�/�8v7^iFC�l��=1�E#���O��o}�)9���~��7�q(I�
��"�0LB\h��+u�Be��@����Ơ��q�G�<�;_`�G9v�~N���͵M�;��ƥ�~KZ��5Z�}D���*�Z=��=�=���`����{�z��}}{�~׸������~����=��?�/��O�;�Ǟ�j�Z��t�U�=uF�����,u�+&��w�K6g׹��/1���Y�$�IO�f؛�xD:�Ө�ƻ��8 mx��D���s�@G���HD8�q쑷�d�ꫨ��#ws��f�y�"wN`}0���n.�a�8zX�
�,�#�п���K��q���A�� "Ɣ�$
�\x��/�C8ͩ�c����$���κ�J���B�ު��z��N�f=��B/�B;�<�T��&K��
�΄g���9�ސ�z$�. �W*�[�g��f� ��L�0�����#n첑�����_{g���w"M����~�w����F#��6�x�cɀYV��B���7���%K�T���e �&�u�Z)�<?�|�r�	��Ƭog����9�0���1W�ֱٌ^ u�����|��p_iKKu�מ���b:�P����(���"ﾛI�023a���U	�μ��?�in+�$ϸ���y�g���H!��I�2�
S�Q���Km�L� /�Hh�����i����7��U��.p��K�ٻNzl}_F� ��d�;��J��p���ˏ����w"ɷ��tOv?��"
�3�y�i�{�)F�?�n�����Ob��,J�y<�:ު#ƶ �'��T�w'���H'.�ɹ/}��7oa2ǻ?�����CƓY1�`9�I��#��� �[���
3E�O��gh	2nWE1c`g\y��o�`;���>��E�\�t�/��0�!�MGxgA��� �-r�K/�!vA).��2��"ٴ`x�	�ÛDQD�#�a�o�}��c����I9��W�ȴf��뤇�(������u���c(��� ��d�o��b�6%�)�yys6����*�QΡuL��x��NA��� �&Qk�(�+��-J$J	
�8\پ)7����+:'�/?����ջ�c" &X��Gy��G���c;���~�����X7E\Ѽ��A���8�8��2����ʸ�t`EI	�t:*	}�"!)��4��%Eȣ-�)A��6'������ed������	�'iH�h,��<�����],���t���C�qU�h��!�cƌD�5~�譗Ho�`8���9W���%޺�x2aC����������cQ��B�Q�V����Y�`�l�{���Z����Г��"�]�̹�"��������ȭÌ�.�>�5.���'��M�>F��
��b9    IDAT��r�u��6`�j��w%��缽�+�J"Q���0��XkI���c~��*)��
)t�;-q0j�n��a;�O����Zr���tO����,�A���{'���P\������W8�}����|���͟q�ԃ����h��`]���&�~θ8|�+�
pʣ���8�]��4�KQ�������f�œ����3Os'�+������h��X�[�X>n��΄��͡V�����n�.��#	��@��j�����y��l&k�^\|�IdY�,�R(p��t�-�W�.�����P^!�~�B�|��د���ף���1~��!c���"͚7l�klE3v�ã���b��lD!��/�^�8��m�W׊���/c����|�9�5JƵ{ʠ[��%�]7�J��˱�A�XٰT�b��Eh�1ֈ�ZUl�2ć�.'�S���'�Igۥ"�R"d�-,I���� �ԇwLh�J3ێ�5O���c�C�-qv���m��
�@��f�slmmA���2�~�K��"�1��5#����(�\�ܥUis{ss;�P����>��M��� D
_���?q�ͷ�.[Uɩ����X�<��y���r�s�&o-��]�x�_�W_|W��1{i�C�(����$�˹���r헿 �S�(i���D$��G��6���/(��em����r������~���f������[���"�Q���;�-�����މ���|��F$y��
��%�G�m�TW�3�XHg�T�.���b�W�,,�e��E�4�?r\�ڒ�Z�ؓ�hM�������ϙ����O?�	>�{�%��] @�ܚ��/���%i��Hf޿�v��  f\+_|�9��׉�'O����G1j��"�ǋ��,ݥ�X�����U���l�B��kʺ���#��[�;;�
Gz�~&i�l�!%�0��![�p�]*_�F��1��c
�-¾V��s���6�[�I�=���<�A ��J.����M��:ݪӟ>��z?��ă�E{渻&�	���xt��=ҹ�ۣ�s4]/�+�\]��K�/�����@���@����o���nOmp�Qa�8��{O�VLR�y�)r��^�cRp��?������Fx��n��낋�3�W�
�*�V�gl�"˅��$c뙊!bc��b� υ�{�C�4��~ѷzư��K�;��3rd�����s���d;L䄽�	�G#���'�:u?.����~�[�}����D2	@�l��Y���5��)�R�x��k2����ܐ[����'PI�ھɥ���s�rH
J��km��o#�.Fz�v�~�Q���^=cJ%I�41eC:�d暱̻�mU�ge��OQ�6"�VLCAp��Q�/	 =L�)�J��Flܾʍo�=��0��8��Gx�g~s�^r�0ٱr��J9������y����Az��@ٜ�;���y�/����m2'8��q衧ٵ[�T�~�_����F����І��э{�+I!�M9��or��W���̧>���w�"�T"̧�H< �
T�W��QL{t��&q�K ���~�"o��e���|��g%����&��R��
�M��4���ź�vx��%[[K�T�m`��%��3��Y�;���������
Q��v��y���A��b�7غ��)j���9�����5.�!;Jn�X����"��`�iiXr����njK������`�Tb�T]��*��B�EhE\RTe0�%�s�˄{�� ��1L$Q��_'.;ͦ5��a���9m��UeռV�HPJ�&��6�au�n�|k>�,3�-�}��d/�ȱa�-�pxl3�6+n�=����rE^̈�;yƝ�C��Oq�c���\�o~�7�����4��N�PJ1HW����*�v�f^����w)%�'�`j2o���,��n��Wo���_Z�{� f˥ힷ������;Ӗ8�m��7���?|���?ev�&������9��O��n2�-i$���"]I�wAs'*�����Z���N�����������|��>�)��C�Ⱦbڃp�Xo}��Kbl�� D��a����a��ŭk!���0��)�8��"쾁��Rh_��*6C�X�u6iH�E쇩����r�e��)D����� '
�|�q ���c��7�S�p���nyoT�a%U�3��)+��&����N��U�S)j�ٮ�(B�9��=�l��;�DPn���	K%�ϧ�����U��f�`.[��N2�%]�
a*9�6��zȁ�9��{��JHF�3���,G�tI��n����o��eĳ�����JU�����-�cGH�`��9������X���Q�>������,�(4�J���({�#Fg1b�n��O�=��3�7�d��Y� s��x���@���r�t,�Z�u& �	��m�r�o}���ɿC[g�'����9��sķo�#�q3���&S�_�h�[/C�ņ_�L�aU��R=���(b�-�T��n�և(��L����5���_=��W��6�[U��4n�l0ĺ�6/�����翄����?�iFO���B3�C��ܚ9��&��}8[��\�"��w��F�QD֟~G{�q^*le]^]T�ҫ�}�y9H_.h�m.c
��b0���m�$��'xwx�̚�]Sٙ��x�-���m�Ӆo��_���r�)�ݹ��u��y1����G�1vY��W��[v]mT�����{�i��@�k8�����$����֐����>�wᏥ�7o��T b������]��
��%׊c�C ]�� )D�F\�<� �3!o<R ��s`A�<��y��>���T�����J����6y�8�6|]��&�mb｝K'�yP�õJ�!=q9P�������s�(Ҡ4Z�,p|��#ڌȿ�x���J��B9�F`�)J��s�!x�D1$�M^��W�7�1Z0�n�2�"�^e��}R� ?Ԥ�M��8���C���g�m"vn����������&�$&SQ<`m8�(�6��k��{}R[WUi��#T�=�d�3G�9ĉ{O�qx�٤�~tⱼ������ҮR�L�	��c�KL]{�>G�WR��!�G$D�%��7~������|���=��'y�s���O���w&h5���I�R�(��~�4RuX���Ȱ���x��������}���F�)B*_��`>M�tਫ਼�����ͣ�%\����]���f�fs�.�{�IN߇!^�u��u��>\�(Mj��k_���|��� n��#��;���y߃l�w��7��������|mB�5]Bk5�K¢�}� ���l��{��+��I�}tD�;��� ��������ǡ�١��D��:Q'�P�>uOHa.ک�&���`K�BE4�ً���Ǟx�e�
������+(�gtڄ���U�^�ʅs�koݜ	q��@��JQ n�������sث׸��_��c���,�M�Q4-~+K[I����0��~�)�س9&/Pӂj�f9L�69��Omn����%����ƣ�D�,ށ�!{^�8"d�j�ޅ(�+<��q�|��﹟��u�/~�[��G�.��F\��9yflD)"Z �>"�J���(՟�����p�����ܺx��[wB�"ݹG��a����j��E����5��X��*B6���*�x�M�6�1�s��-�t�7��/�/�L~s̱'��=���m0q��Q��~�^)�v-��.�"KF����a�L>Ef7x�+���6����Sl��8-�J��J�[j/+"�qo�s�,�}g�ΙSlڂ?�	���_�N��ɩ�A'X/06̩���BT��_��p�x�+�\�<C ����I�²1��^���7��>u���O��鄘3�����������uF_�H>�R�Ei�s!Y�m��=���~�ZB��b%�ύVj���w��*5��o��bl[�W�T�몗�ή�|}����]���8�_��4*IpiB�������c��%67L�c��������R�:�N������i�{�H�``��<��A���T
��7q7o2���|d��6���w}S�k�/2�@��1	 �P������,VE��67^���=��#�YA����R��YH�4��.Q��Z�}�~�ͳ�Q�Mf���op���O<���7��#���d��L�s�6^��u�.�ܫ�O��]R��#Ak�f2dd%����I Tj�|�u�����5K�#��Q�B��}WG�]Ｊ�ߙ��J��!� �ӽ1�T���������9a�+�}�r���fbU�?�w�����b>�N���h v���6��ˈ�ap�nN�c�#�VeJ�p��J�����Jk�U�D�z?�@a9���=vo^G`,5ɑ�Ἒ�^��o�U�Tg��;uƱ[��fd=u��1Γj��Kor���wI�F��x�pem¥�5iF�aZ���x�o��gEpo���]���)��#�2�<XH���HF��t�"�4M�{^ |P~k��HC(�PA%#Ps�ĶhLC�!cQ��:$-\�
�A�i��x�!C�R�!,�<]D!c�\��&��^� @���'@"��eDC�s��E����ч�_�����G���HH�SQ`��XA�$���<�q�S���\�	��q�uFi�F'�x�*\�� ��X�Q&�H�є�%�I���������1���J�s%��(!1!�Y���̿��CZ���k�k�>�g��m-�b��hw��s=��8!W3.&�����c"��s�/}��J#&�0ÒF����2^�"s��_6�$9x�pGZ�T�C$�鐋w��}g��O�;��/��K?�!Z;�l�aD�@>�P�6��X H��!Ŧ�xi����L����(�f&3`�� ����E���W� 4|�=`C��=3�F�"�(�p�Σ�Q��A��!�9l��V�-��I�#,FX	K��T��q��^��(��@%�u��Q��V�|�*r4�L��x���ZQ�R^&Q��<'x��~���
Bx�O���&��1&�D��L	2� \�pq�sW�$wx�W(#�t%zPB�n�ǎ!���˯�9;��3N�9|��O�ͭ�%4�\c��=��#��}�R�*�\�3�6T��^�4F1����I����rm������v
w�I6�9����:�$���|�W1�(k�B-��"l^*b���i҃���ք(5���W��+/��#���&�^��df���il�AVL!�a2x�ؽQx\r�W�J���ґ�+	Zέ��,iA���h�%�B�
��I��� �>����!ǀ�$)Q��f�<��[�t�9��"h�|e��J�W�!��"�q�����>(�����_V�sdTI��E�ǕvI����/��ԈB݂�Ug�w-�zu�ȶ���_߇S)�pH/�:�(�X�D��1+J)t#TDQ�1�#���5�u��M��T�B�F*�����ǚ�2t�0:�ة3<��Sl�P��0�p��
���a�F�����6�{��UE�õ"s9&�!,�rꁇ�؝l�s��K�^����H��Q���3�^"�g-a�'R��:{�#}�A>��_���S�1���_�k�l�u=X�4���ۛqaS+�92�)��0�1��ʉb�y�~Pɿ!)Vhk~�i��\o�V�%��`!~[AQI��Uuj�W_���#e� �Ϭ{C�G�0�`K�4�j��rm��k���[�S�KWx�_E��G����{���1�ͣ%2E����"���՚A �BP+�f6!�y���+�)���Ü�Я��:�n1��)�T�x�l<Ca��l��Jr���a��{����kI�\~���^�8y������(�y��^H~.�����u�U�����(F	�@�DN0��Ę�ȗ��tJ"#�Lc�5D�H���������RJ���i�Ь7���6���㝎9���j�4p�X�_}ʃ�z�7T��]mP���w�T]P��ڄ�>�U���	2����5�wdɀ�=���	
�0&�0���2W{�O�c��#��U<NϢ�JbT�h� ��,r�8j��	W��~����G��U1�h�[[��6�;��~0^U��D�'�$���܀c=Α�ũ=�c��96�c2
�v��^c�%�ed�c�C��M�w�l�ru����r�ϒk�.p`��`6&���f�1��X���"����H�0yA6��*&Mc�0HY ʀ6}Ġ�}A��SbS�D�?�zV�N�WK_[8-\��T�6����(�e��)Z*ֆ�DQBf-f��_����^���oD���\��W����`���D��e�D�Q�@	��x��.D�,����9���l���O���շ�i���8�}g�)�0h<��ܡE�;���eW9�꼂�;Z�h�yƕs/r�G?d|�����C�sK�<*�qX�a]�	}n��S�L�X�}�6�gd��������"��~���yw0�t'd���^�D9�v&��c�Lp73�K����/�3�+������aT��UD~A���.h²��v?7 ������R}��@�|���d�:�e�ߢ�^���6TW�i�C�X�"�1�d�Q�<���"��@I�t�to� �"�����2�Y����,��Z��U�9��&R��7�!B>�83�8cv�"����h�B�|����ݑ�l�o�v[�x�w-��)(lN��l��N2��Hin��2���10�|b�3��,Y��9ܪ�X(
鉣��y��IG�sɡ��r��>��,�O���/�ĥo�#Q��g��+а�M炭�d�I�X뙭�߈�:
�ٙ�[O��ɠ���:�����O� Ј���O�k���m�_����7WI�#)S��Q�p!��L�%Y�D	�Q���gB:2?���_X�5mx�ā��]��|��������8���2�8�N.'3S�R���+�}�EB�,�$�f��~�~��=uu�F�D��c�8BF��zw0�f4���'�w��UOaBIt��l�hz��8BDd�5��&cJ!��8R4c���6�_%അ�:c��88O���cI~��~�sf;{�����~�5�TX������r���~4�x�.{�u�Sj�Uˠ������[�.=-SM��,���!�r�P����k��U��\��W�^��3�:��,��{1��4�`��}0.2R	~ga2��D*�9Gn�F��2�/ݿj�<�V���V��j�ԸC-�Ŭ��cZ�S�?�$X�!f{����,��g3��T7�oU��|a���~��Ǩ5�	�oe�0���wq����S�}�W��-��YO��J�3�r���\�6d�a.�@�<ϑf�Ipm���Ȅ��$�<����u.~�;�M'��%I��iI�-�H8_���O`l�R���+��β�Sn%��m���U�����ZյHC���p�!��CHSF� r�AH3��Q������0��(��ˋʐ+��ȧFD�x�m��#L�������8�:]��ud�˖?K&�9�����R��-^�ǿ�\��^[��G>�ُ~�b�0�VH�GQ�G5l�U"d���`C"A\��������z�$��;?骎���t�L�1�0 � A��YJ�6$qcC|R�bc�u���Pl(Vk�Ii)�A��0��oo�ǔI�YU�N�:�6HnvT�����������:����<�U6N�%�#%J�����ݥ�}{�gm}�a�w�=.��c4c-��|����9.>�<N�x�H�-V�g�9딪�y���m�|��s��JL"p{׹��O�wva��0��AI"�ԍ .|@u<�널�y����W���{DZ�^�bA��ߚ{#����u�N�X�a���o������ꇄ�4�NjM�b���Q�]��r�iJ_C��%��d�[�3��|X���D��FXa�Dg{�~��fx�(�!tģ�!,����#��k�;��v�>�XĆVhbx���Ïq����3�7����\��8�    IDAT+-F&c��ͷ�|�-I��"�roA3&�IM�P�>0�x��ș'g,�۟1��mt�㼊��E$�R�R�V5�@�%H(�x﹝����\x��p���?f��[�>�w
����;�y����h�&
�	C&Ӏ��<������9��/�'�ԝu�K�V�<Tվ:H`��6s��O�S�j��D���B�1o7}1KV�'mA@J�֚a���W�w�~�_c���\m��[v�t!��<��Y�K��19`��,���R|�&~r��Θ���k�ؕ��T�����{Hs���Q��%Gb'����x���SO����Oq�9t�HS�D������~�}�{�AV	c�{�����>x����%&{S�>��z�K�jݠm{03?�q.~�����u�Fxk�bi��B��;er�Sd	�;-)� /le���-JBي/��m����m�Ro����U�׌�B�Jd��f�}|�^�;��^�L���v��J4ldbre�Ir!�����`�ô��s��к�t%���ޡ������ii�B���&�~�O^�)�����Be�Ҝ��TĦ�K��m���%���8�2(
A���g�"7�̲;ȫ7���L���e4�yق�]G�ݶҷ{d����GZȝ'����S�B���u>��������r/!�x;ŕs�b���J�R!�N�0;�f@���s�Γgw��e����2��7�E�"B��8kK��Ih�KJ,^D*�CBq�~N|��x�����ɯr���q�2j��k}�ty���d+�C��X!��a����k�z�2XK�v�ߵ��)UUf���i�����o�/�+/����ӿ��L��bόc4zK3�[7]Y��v��MH�
M�5��%7^�	[2�=Kr�s�kC�y���Z�a2�a� R�xQ���[�~�&�sm�z�Y�#Ǚ�bU8!��9�g���8-�c��& ����^1����5n~�>))��M���R����W,������=ڭ�ƅ�w���Ԉ2@��b:'����A0��1NH���B����r�p�U�M������A7���n�B#8��[��d�y!��(�("���{9��-cE$�v�SJ-����51�BS$�v�ﾴ>�LW�i��s�5B@Y�ڰ1� ����׹��$SS��JJk+-h!l4����[<��pl����C��J�Ԋ2V�nn�8����ĵ�>�}Q:�,� �a/Co�n�gH�_X���y@)�
�%&`vv�<���]�;�x��ELw$)s+@jD���b8�Z
����@jf�_EY����;w������9��6�_̙�BaI�]w�l=õ�x���� �Ђ����7����/IN�b>�P�Z����w}�{�#��h��&�@0_�x�������r���W�U��1�_��"�ʆV&���V$�b����bb��x���[�;Ͼ���m��ak&ҮV�Q��˷R
!1�R)Lȹ���L_��r�>��Ϟ!M�(!���D=��N�4��3ʬ@(E�Ǩ��Md9�X3K��UN?�89%E>C�V����1��q�>b��w��TK�pR�0����mL�(
/H�!�yּ��$+��Y�i��RsH���-�3Kb:�L7�MN�>��c�р�%^	�
�T���E��<a]����8]�]���ݬ�6��A�N��׽�n��kZ��d����ϵ�C���DX�>��M�k������`��P(��h�AH��4%�#�T�a�-��&� �z�q�T��|@i��ǼQg�[��є���:���#s���;�rN��1��	�)�!��-��-F�!E���d��RvDdX:�d,��|@�z�� � 	D�HP�"R�\B�"�=HO4�W�y�47W�#V0����,�6����O_A_���Jq��!�܀T(�Ϛȁ�E�x� ĺ��h QB��zΩ�SB4��`�@di(���v�y�[�I�a��I殰�MI�cv˂a��}$c�O�~�)����~0E�U3G1��dꎲ��י����O���wAc��˒��C��bci�I)A-� ��"����m)81<��t��/�����a��f�ὗ��wC�=E.b b��Q�`�{�hT�L�1(�Ρ�Ya��u���%b}�%�r�U��O�@>���� ���)�I��y��� 6� ؼ� +RVu�Z��Pa��K��ȧ����Gĵw��	��M�g��?��Zñ�a3sX	�p�0�tٸ�$X��� 8�A�}�(�[�[�Nl�G\}���m������q�/rEiv�g0�QCf��`� Ʌ%��'n�lE�$����;�s�e1)rx��8�0#MA�,܇m��fu0�se�P���AJO��ݶ��d�
�Rbf��(�Kfh����f��0e��3_d���k�x3&Iv(�	�*ȫ>DG�oec�>/���@L��Z��D@ƺ"A��[N�q.��T)��!G��=d|"'�7�#�:�0��%��R�֠�)��@�y�t�b$��+��-���q�D)��	ZF�
U�<����@J�(J)"Р��8�P�P*+!���sD��	�h]	�>�=�P�:"+�`E�ģm�KJR�J���5ٳPm��V���D�Nk���0�յv���ܧ���B�ƚ��g-��ɀ,˘�S��H-�;��S�����*�(�k���zq,�i̻5z�X>*���D�Ek���{iW(��&�JD: ���֢M��6�x�;���:B�g�i��!v�`L�#eD�2*eg�$=�4��tF���yN(m���eڮ�Nb�P�����'y����ęS�^����1�rY(�0J`�m"w�$��5�5���x��*04C)ߞ1lq��O�>p���M^���c��Wi��V�T%#i���(P��\]���R�˶i�~7+.={���o��;�q�\Z�봶�bS��������S�N��ڲ}�_����=v�OO6T�Cb���b>�X�dB �l [CY����^������1eN���O����9�Ԕ�}\�a;�|�9"��sU����%��o�������;3��ǜ>�|��[N�B�ʃ���aֻ�����U��$IH�F��>i�z�6A�?u����C)I"4���~Fz-m�Y�:t���q�Uø�,dd=P7�p�ǯv���m�s��h��d6���QHuX�Y�5�]��ig��S��!�Bm]����As�ݛ�9�*|�z��ܤ���k�S6y�s��k�{w"���3/-u��y}�f�C�;ˋ�۷���Xځ��#M�Q���jT� w�8��c���˦���c��ݬI�H�c��-�p��#z,� ��[}oD5s�3g��(I*5s��G�8I��8�ݽ��z�.Zr�-�Y���LD]"����;k�QT���<oN���^��`�I>�1��}������C�����a�6�QQY���s����9�ŋ`<��~��/��E� �Yt*dDm\1�u���l� �h3d���g�����G�1-���\��?'��91�H�~�{Tr�V��MQ�Hc�!$�S
� �X���6��]���f�r�_\�o`M!,�b��U��d��5Ԥv���G|��������J����o~��G����Ҕ�,�S�6�!Y6�m� PV)ODk�􎑑��.W~�C�K��P�}��G�ǩ���`�,о�'�|�H)�P�I �����з��bș/~��'!���]�~�����������{2΍���9ʛ��{�&�Ol����|Dz�)�H?��)mf�.��=�>o(s_0K���p�������3J,�dHY���2��F����f��`���?��J)� �C��E�2���ǧ���*�j���}�n��;4e�z�5é����Y�#�=Ob< "���Y�C���>�sP����E쁁�e֑9�O>I�Z��%�I�J���Md���ih1B�9cQ�n3m/���7��+{�O'"?8O@PŃ_z����0�\1A���W%5�Xd��+ʘ=�y7������w����/$��Q�!���I��%av��ｇ��RB��_豴F�@��Qc6�?�C��v��c��d��1L�%���r����XK Oa3����;�6|�p�W~��AN������+�n�`,S��$�����`�?��n�R!��tw��A�m�[�����C-l��������H_�uh������nv�k��d/����.J�����y���3ӛ8�H�)s����ĭ]W��������&�M�ѷ�����-Jf�c�<��d��iLmꉦU���6�K�c%(��?A�!G.~�?B�������1|�~Z�
��7�5R�{7���Op�� ��i��0h�Rd�����_�pb�?�� }������n�"���i+ <���iK?*^��R���:,_�ފ�����S[�,��ݹ���m5w���mP����~��t�=j�t�Knb!�4��Π�ڝ�vk��D�mί�i��!�,rc���Xk
G��.Ǘ�a̋�>�y.�ƔB���R�T�Z=�y��&_��{A��iw�v3�RؒR��.�C�7�!��7�S���t��J��L�d%enu~C��2"�:��^_n黅��9Ǥ�IN���_���1:����bJ"*�6�qu��)B��v������׾F�|�^"�3�3� -#�
!V�+]3���E�|:����ǜ|��x�[�̝���q���Wy�������-�I(,��[k�q��N,�T�RJ��Yg��(���U��A�F�^�:�P��F�:�}�.ϸ��"6��.��o������ٔ������G�}��b��F2��"�rp�]�Mi���<BJJ瘗��$��Ə�=�G&���|�����zQ��`8��t�}̨���ZG%�,&���g|��+��Qd��-�$��k�1��� Z*�C�J,��5�e�#��b�8�y�w���c��|�n�����5��=��C?@����t@���>��*vD�]��`E �!�C+�r��V�J�(�{�|fitǻ��ْ0Q׺��dr����ܓ5�$$i���R���.a�����S�v��(˺��'��e$Ū��m
-��:�B@%E���1�ӈd�3,I�1�u����V��H��}�a�`�8�x�﯊^�U�_���]J=�S �S�"j^j4�H� IAq�2�(P�&��߷�̋X,�)�Ojm���X
�qcwa�\�B��n�FtF�M� غx�����ѐ��en��C݊_���X&}k�M<=%�N�b5��|�٤��O~Ļ�}��X,�$Z
����k�
���gcs�������<�c��u�.�g�J�_��������li�������a�5#�ZSzGVx��䮤�!h����jT]V��nV�2������`���l�O�'���CMy���q�����o�-���}������sub�A�#5#�V���YM& '<�� �&T ����v�}�ro�p�8�|��̷��iE�M�{�.!��\��%Zj��y����\��a��m �>Er�~r/p~~���?��ۿ�(��"�v�%ER��&�;W@Hv�~�SO�@n�Z���F�g�[���흃���;Z�h4��hu�<��s}?����ٴ�zI��ൾ{���N�[��A����^����t��m���ճ��|��&��
�!���Ж�]_�A�c�}i:X�,��e??��&i��^��b�$.��g%�(L:�C	�=ʽ;�R�h4���j���zBҷ�Ѕ'�Li�գ��ʂ���h��!^k����ϥW~L��"`FY"\�sK-PR��ti��Ϻ���vm�Qk�AD�TP�%�i�
�;X=��ϸ��|��0���@$*β�C6~��}�&��Ǟx��>.g�w����b;6����^x��R~�,A���;�};ESf�g�ǜ|�Kl>�(�+��2y�\}���?��|��)Rl4�+j5V,!�F��Fh�u&E��	O���[�;��wJ|��T���Ž��=�}�#�'.C͆�B���On���+\��f��w��?�y.~����9ؤK�8���ʸ����h
mi��.}�'/}�d�Ji�.N�e?j�<�]IB���/YybE1b��:vRI�y�٥�щ���p���ǢX._���?�:_7�J���V�N�
��܍�|���b��l��0��b`��E���x]����a}���3W��p8J���
��a2!
�?���9&"��;P� ,��u�T����6�U߹��P�(|}�o�ƌ��kd�OP����m2v0���f��A�~ͩ����� �~��VM*���[��^Z���/�*�1H)1j@�9r��h�Fb����\��#lsns[��y��B�op���^�W`V}�u�~X5�����y����NI�`r�&��+hb �oR��A�27�v�B��w������J꒝JQV�B�G�Q8����]����#�2��� Ix�0yn��<��W8����"�ꛯs��W��)a�
�pi=�t�h4�X��Ԍ{d�+���{���|���/������ǆ�Ǆ0���F1�4�i4�E�B �$I���mQ�"�|�I�"��z�ᶠ���u�{��H��)�m���=�L'B�ؑBLJB�Ē�psr�r0�����?��d�L�<���x�_�0C���\�^�})0J���!,x�w�Rr�w�\��,��N������6�|e��9�Zb���j���j� ŉ��0�|��~�2���:��yҔ��*@�c��h�J*18��U�R�0�e~���2�w����y�\�P!�I��=���4��~��x��_�P0�s�r�bF������pw���"����ג�,>��HŊ寫��j�-��:���k}��t�o�����6O���M�F�Te8#4�GJ��Y�
�*?Y�=��B�@ ��*2&U�Q������"�ȅ���"�R*������$��Q�D"t�:�3 �BJ����"H��>���(�D����q�˚.�߽�-��Wp�s�&�A��쥟���ƒB
FN�m<6d�S��b���
��"�B���j�4�\M��.4y�h�r�g)���+��`�^=��w�e�<r[��ȡd�_c�2��M$�
pH�(mV��h�(��m�l�Rl��s��ޮ�`2RE,ZIR�b�N=�􃏱u�n�9�ܣ�{��QJ�L�S�rW��2�R���M�Z����^"(xJD�)���d�h�4���$��$��'�����.��f�5"H�W�4a��,gCD�@X�2�U
�4>@i�v�A�m2u�_d�s�����|��~�?!߾E�,�p�JRr�:C�(��YRmH���%���=����Y6��>oQnJ�K�Q8Pz�P�ҫ�uH
�V1��v��@M�q�T"]��+�Q"6�,���A{Ű����ܗ�D�he�W��e�zI	�;�����=e�H�*<[�����v�Ý���i�c�e�+g$Y�N�\dO@V�"��8� 4����a��ܳ"9��q��O�'��)��8�M`w|��dW8�Ԅ �֑(I�%��+�B�F���R��#�!��&���$-�dh6�1ߧ��\V�DF<f�T��; F]��VX��-��1����dR
��,L)�"�RϦ���	����8p�l��<���ZA)��AYх$��E��d��.��V�}n)Z����H`|ms���?���-� �{��ws�x�D:�הJ�"��꺷?;B�g4��Tq��#�!("\zPiB#��Uf�GV|."Jh���U�7��&�b>��q}T8)13�R|k�{e��B��@+��=b`0B#\���d�E�Uɼ�s/Gw���.��s�徇����h�d��?K)�b4��&MS�N D� !,���;ѫ���bR��K=w�z�������7Ʌ"'�˂a�Ѕ���~���gi瘪N�j��ޔ�t�0/rL�R��t�p��y�,��I�    IDAT=�(�z��l�x �߸�P:���l�?�N�̢X�̤"٢���rF�#���<g�5(FJ�e�ظx��>���QŔ��������ɋ��U�{4�sXׁ��֒�9d)3�r[���)"����E�V;o�1�k����m{���.b��u`>���A�P	�
�����E[K�/���_�?�?���.�4�ع�9��s��-
UR�%޺��;0��p������7~����X'�>Ϲ'�g"v�QS��9GĸP+4�۔�tBZX�|FP�m3x�4�e�k1;�ʹ�]�>�}�Nˬ߹Ԋ��cnOf��%��1�����:����{��Ż�J��cq!��|�%j`H7��Db�HZ��kW}���_7o�������.F��u]�������:˰se� �葉�9A�7�67l��՟�G{��^�a���#ۻ�5�t��.Cꛜ���'�A �&M�hm✕��RV~��0׍�o�����6���xa%�^�V	���t���I��e Y�-1z-��0��1]#�����:#�4L�k�؛O�~�*y�a��ٹ��"/g�?����fXi�}�4��\h�G�DA���3�=ǩ�!�����>�ĶR1Eh���k�=��i���a�H�\��W9���$�"n_�x���	B�
/!jl�E�\$��쪟�E�N���JnKd^ ��D�Րm�2�00 G�w���]WA+� \,;���y���G���Ec�l�s�����mrB�8�����|���-��y��_�E��#�U�z�Ui;u�N��C��wSF2���b�:����\���ak��LU��!�� K�fkk�P�sF��{�ٕ���1�p���z�L %@ڿ������\��ꮹ�q��}J�}f���%OQd�)�zA���+W�R�.�����R�dG�術��+�h����҅�*2z�txb`��S:[��cu���~�meQ4�hRʕT��o�� O�=���-}�}W���A�v����Y(/Rj��|�mf��t������Lb�����m\�E.�2Aj��>�L@��t?ǀ�LP!��	g��d1}��Z.!���t��W��ۚT)�;�y'�2w��6�}��!M'S\V,��;�Yw>z~��`;uk�ag�5��I�S*��!G�?�3�=��O<Ά1�̑nn3�������1�z#$Ey�����s}�=O!Gy�ϳq�(��y�/���ǟ�
��6ź5���/>�����j/<�sG�}�SO>�L@>���������q���HM"�+�/P4� J/�%J)Bq��4�:��r��x7Ż���bxػ�j{}m�+���$��-��X�`�N̔i"U̾'�y�(_0�{�7���_�DF����l<�(S%�F'����c�� ?��\Ok3��{�D����"�(Ԉ�3�	�`Ii�i���ޖ���s����)�;�>������.f�'�2��Pj�kau�������ٗ�T*�x����9~�!N~�I��9�0!5�1}�d�������ںiQ�B/+W2Tk��Y��>���EU��y	O�A��Z�r���w����FL�^��'�)!��1Ƨ�察e�]2I��t_�)�g�[�/~�3�$�&ǺÈ���1�F ��5�,%yWFM:�4�5&�N?�����PT���[��h�m��l�t
�}��=�̕XW���I�hL��|��	�{�w��߻��Q�,�eI �|��D ����x��>�h4b��.�._��'S��1H�,�֊�� �9J�ذ!�'��s��L��Zt���GOP��]���*�f$���e����ɽg���;��'>�%��y��wnp��1)'X/[P�� �\�_� !%Jk6�	��j�ޑ\���RjȂf�'k1��v/��9������>��A%\�pK���H��h��Ϫ�j	L"[���|5�R[��v��&w��}��/~���f��^�Wd�N+���KD=�{A�{�~�׈�h)� ����@i>P�r���Q��0� "��`@�w�[ｍ����p�$�V�R+�saFj8����{��n��߭/�����>�ͫ�����s��3c�\�[����M?Z��1�uL��� 	A�bL^��� �
�F����h�/ �ˣ�3���>{�_m{_�Z�-����[i�3����K�޾��7x�w�" ˼��6y�S}��?�%�]���Hl��>��_�.��Z���kYp�U%	V���w���(�����=�{߀��p/s�(���V-� B�%4V�`HQl$9�'�V��ܦ-��|�G�|b�kM����>�$᳏>�W^��w���ի���ź�t�0H�$c����໨T�G�k�Z� |��Gℤ�'4s��Ot>%ѱ���M|X�t5�o��>�޻GRZϑ��7	��0��ob�n!�	$�W�ߢN�Ԃ.���hV�����w��O������?����S��S�Ze��t��>m�nG�[�Y�n!8���s�W��GNrm. ��P��5h�H��j��f�V����6C�����v'@���}�	0�.���R�0Q��"�.v�n6(\�����1��Gh_ �[��Nkr�_[��)�r�R�E'�� ��9[ڀ���U p�����4����ۺ��������]���#D6Ë�y=���F�;�η�����X �h��J�TY;u�,�#<1��� w.BWkRc{��{��Ϫ�*�n�u��}�D�%kj�-�"
˫�����=�� @D�5J9�'��@I%��,	)!L�.�?��t6ԃ\.pP�.�����w��7!�?PV�_�c�N�QW�DU�Mp�f,�_�!��D��D,�")P��Ɩ���Pf�_�D�O�|�M�����};HKl׮���oIJ����	W������lʄc��l�҄�9Fmn!�����q���Q�+}j��+�A�*78u�4ag�~6A���e̊��h��ځmB�X��X�Sngt�~n�	��������ݿ�q�ܛ�@�z׵�E��}~m<z�N���_����.���ȗ�����昫���x��۝��ˮ� V߫ġ�!��W~���Ϳ����l��>��:ƥF�l�Pi�]Сv_%�D%��&x.�����C�)vv���/�6�x+�*��+!][�Z�vŌT�l���K?�!���l��?�pg�·��7~캚�����b@�+-Ӽ@�Ău�rp�-��+�Y]]�k���_}f�uB[����g2�p��w�9J&6����D+�h8<T������,B@�'�ʪ�*���%��L]�����m
)�u}_�_�[}���m�r����@����9-X]!��������כ��=W�+K��{;�����^�횉�Ei3ضo��ݏ�.�}~���_�ׅ�)��ٶJNV���,
ݱ�C���T�@��{s�#|`s{�$I%)��_����h�}7���8����u�Yp-F���#���.c�Iܢ����]��;��@�,�!R�$��Q�k�,,s�'��E��׿��sg	Zr��gX�#L����dw�	2@�$P8rk=`SMy�fﾅ+�H
K^V\^t߷�ݰ����F�_�џ�<� H�&�{w����>�(Ѻ�꾫���^'��"���X�안�S<�����+�߷��<� P]7J�r?�x�$#����8��{�Q���vN�г/�q�(f<�W@U�tZ��l�&h���9�l��e����������O��.>����ft+�a���u��B[;�͸ލ�{K�gxe�9w���?���n<�a{� ��ǐڭo?�i�RJ�	~2�Oge�f��[.������Gi���+�.k"��qe�-�|�8~��ΟE�R��X뱅ède�梫��U��������v�ƿՂo�3V�ӟ��}�}�	2����FR�{��� �`ʮ
rX�6P:�:�@=�
�"���"qx%:"���#58��3�!��G�*��BE	[�X�^�oI�n�%�dE�㘜��;/|^5�G}�'x�u�dC��=��� ���v�C�U�w�
�,sUI	"�C��dD�
���k��9�Kuz�\���ʞwoA�Ҡ5吉(�>q{|�K&��W^�	�� �T��n	X�5���������uO��R-��BA��v���Pr[r�0v��K��~�~�l;E�2w��1'1n����� ���2�!0BRj�P9�� �D��4��S��^�����.#a ��e�`�9�i���d,8S��p�b��g�Y�'_�_�wt�}�����z�cN�e�` ���U	��5L�B!��(�<�Ch�0�&d�g�H��9��
'��cs���Wx�����ΊM�Y�JRP����K��"Ȁ�����"-6�
?Cct
R₈�C(���XMH��������}�(6�}��~�_p��ܵ��$C�H���<#����`��vU[����ۜL���W��|�-�,C�?���#���9j�8�'��h\у�"�ZJL��Sl'�b���>�tJ�~ã6Ƙ|�(�칀)�S8��k���ItP(/	l.�Dl�:��[�l���gƈ�K�I��nJ�����Aļi���̈
����
�[6n�g7F�a�a	3#��D��]HGr�;�-�p�w�M5ʗ�Ļ�akQ�)��F!���T�z���:�o�s7��	ň�X�W�M�	lL����_A_����Cl>�"�/�	�V3���M�|�2i�#��j\%�ǌ��\�;�8,�+"������"ӶnJl)�V<
�" dB���5�
�u�Ʋ�8\ۅ�o�E�.z����=B�:G�%e��T�0
4>&� �cI[B@K����-�蘦�����;�E&Qko=)���v�#I!��~�u�.=�-5U0�"��/nm)��uM@J�X	b�w�s�}�ο
�0A��Ã��O��EE0�k��6��f�{��u� KL��,�Uߏ7woE�	sSwm��{��6GN�A�	�@>ۥ�ܥte�x��8�{�ΛW��x�V� %��l١t׮]������ah�ͮך�1�!I��Z�p��\|�)6��+W���7���,"pF��nYi9v�8�K�����[�c�ϒmJ6����~���['��Y��e��v�h��r����+<J� �HH�Y\�Ʌgc�����k�g��s�����s.~��월R�l��
d]I�X�t׎�c����|��%ds4�,w�'��r�x��+f�)�9L�����KOń�s�
��b EV�t�0�bA�|�ay>��g�JJ�('�&\����]�2��$*#�c�"Z����F%+�r��v��Zf�~o�k�ⶵn(��1����e�L��D�U�om>P&}sҧ��}iO|V�(.��(�)�o^c>�!D$I)%eYRι��ܧՅn_�ͱ#➴[�|�5V!JjK�j[;�׭���v��a�;�4�5�9m�w��i�|N��'iB}��)��<�܅ ��^���CG �;�Q�}׶�#�!C堗!�9\1�����꠼:�(�:~�A�<tJw.��T&�#Z5��Z�D(	�w��@x?f���S�����:%�-0�����y�x�/r�G�[�̕��#�NQj�2�y�MQ2P�XX&��@�z��M���W(�B�H���M�h��%����Ŝ��*��
�X�+�_�0E�����I�0ۛq��w��'/�-$&�(#�#r����f4H��N���l~�󈡧��u�|����lF��!;����ʁ_%�-��:һq�G�-�ڃE-j�p�^�36��!��������_v���n���_�gy�r�#�&�J!1=�~_�H�6�/,1=�t$�d�����\�ǜ|�E��-%y�B�ʹFh�c2��6j�>�|�t9r6A��>v�앞YQ��A��ф�k�k�

%0R1�˸����.r���a���d�;G"UcMjӁØv��A֋5�Lw�Hr�=�v�������IY�7�G�ۊ%����󽶾k��G�Q�l���M�H�0HG�6
�T1���0��}v�Na��ܚGAQ���+\{l�XXz���
^�^!�&�V��s?�]���e�N�}�r]�ߝ�����b�]�S�y1�������|M��L�ҳD���Q���.�l�ͮ�P�ڬ�J��Dm��l}Ԁ7}�G8a� ũ�z�X���h���d R!���3�-#���-$�.�n��nVC����:�ar�����W�|Fb��y���݇U
�l���N�r�71�	CSU�
r�ɷ[#TV�ƻ�bZ����H-��a�G	�@��)�]��BQ�'V�BȄ)�0:B!c
��}{�#	�z��Į���7�2��l�@���Γ���<�4[�;�k�y�������`dȊ�b2C�fK̽o�t-,��ki�B�җ���!H��	�t�lZ�a�;Wy���+/��i�Ȏ����_⮅4M���FI�X�,�
�E�HT��Dy;��;o�w�
&p��'8��x��&�
fW�KOq��.�9D����K\�ǭ��#�~�A����9�`�l�7?!Dk���=;M�XD�V�2��]�$�J�(E QI�K������D��\��s�:����]�' �gZXPW��
Ǳsr��g`�0�sYe��i�Rj�v�!�S�{�}�rQ�iq�ų*-W�r(+�_�Rϫk�8皌�z��5�1����_�I�@̨P��9bx
�����s�=+�JK�Y�?�&�?��>���D��������Cn_[_���V�[����:6����׾���W����*�#�u(-���!Kc󫮄�D�0� ���b�5�o3��wJ���	"�u��*���*Ӥh��	��$0T9� ��`3U	���ɷ�>��t�`{��ZP�ItQ�����'q����v�=s��Q�T$J2�}��^y�?!���T������a���\N�D�}_�b���fs�,�,]5�Ք���/c,@���!�(��`��̰��;J�"���������)(�%�dN⏜�_�5����9ӗ^b�G��@Iz|��
a�u�F;��W���J U UB@�}�1�(@�C@%G�*-�Q���'|�_��y�\�<��]�a8E Wzd�K�p$�X�)z��\{�u.��6�9��w�?���W�$������̪��m�z��{zzf�!gH��H��!S�˂ ��?�?�˰%@HK��$�
�Y؜����o���23"�8�YYYY���� �[Kf�z��=k� ��S*�9��VW;/%Z^�ޅfs[��������?����=����ǫo�Mr�P4�C�:������H����RR�P9���w�{!�`X�j� m9��^F����V.����˃�kG�q��r���
���6�&�?=��2��Q�z�2Z���}�� <��pv��֫�S�x�lO9ҧ2��kޅ��E�=7��d��*����r)ݡ6,��0 4���3F��	SzN�;���fN:=���)1�7(�s�sv���3� p�"0in�����}&��w�3�m��L��9������Ԗ�)�ÐUV8��IDEѪb(�K.HN��|S=X7�%ȋ$�!g�r����J�*υ�����S����R�;�ϸ��#֓�m���9�*�U��B���ʊ9�]�7ׂo��4L�~i^20dE�2�������-^��o��-��	��h�@t�+������|nsT\��h�����.����x�7y������O>%Da�t��D��k��[��i�$�7�(��C9La�4tWV!�[��Rb��q���­��Η�����H<~S!bۑ�<hR����g�-�s&J�	��)��?�v�
�~���9�s��	��"�{�!jm�[���A�UTU��+W�|��g��Zq������*��*XA+E=T컙�����Ͼm4�#\�y��k�b���q���/jK�u�O�*< ut���O�ٱW!�*\�-(�#�ix�Ppe������0sS��Us�q��&��~[�����1�?qZ��y)�    IDAT#�Wc:X/f�9���7�`���0�;�ܻ�p*�����I��<�oN�q&�蜆6�Ԇڌ}��P�Ԗ��#B� q9�8e����)<�t�G͹��.
x[��ܓ��� ��u�'�v�<����KD��ܗch|:���9V��N xrI`}�G=��O��9�s��?��]U���w"$q��Z�x�}d�o���Q���Ჲ�j�d���b�X��o5��#R��R�	�%H@��[�*M�F�'�'	��`_� bN)��]y흯����N%䧏�>fUhb���۫��`h밢��8�p���&���l�\�Җ��}v�~Ȧj����mF�.��S���M�D�PCc(��,�LF,<�D�'�t�٬jv�S��A�m[�}�	������g)��_G��e�*��uE^��|�#�
�8!;O]6��ὢ���}:h5�:%���"&�f���,H��P	T}G�9��BG��X���v����pIٸꀳ�%�k�����o��U$����꠸�F-	K{妿��s�xʼ^_��W�y��b���*V2AN��_=X��k�2V���H�RSD��pq�
،YT�*�j�)�����Cf��t�4�<F������QL�|�s��艹<��VT�c��%&30�s�� �-��X9�nل1�r&�(� 9.J�G��H��T8��?3yF��<%�4QFӸ�!�gn*�̙<�D��Φ�V>�j�C�Tg�'<F�0K� !�	"����׋�|O�'献�k�l��W$�\5�~�V��NU��]�ԡ�a/�9Y�)yq�+{H�#�$�j�C�ێ�����И�H��('{b:�a+HƇ�j�B�q��}v��9��)O>���ϟ����n�*T��a>/����F��zV�����w�������_r���w-�:T*�ړsd�=�$�-@K����m�PE�t�X��Q�Q��7dQ�U���Td�[ڔy��O`Ms���/�Ʒ~���D�4�Y��A(��=�>qUMĪ�iۑv;��+�1��[_���͚�E �T�Q��Z��H���M��{�͊>e"�쵒�]��UA[:�}��t���	t�!}��� 5]]�o~�XO�����ĺ2osz��^�a-�Q;Ue�����?�.��T5����;�@���`����u�C��s�y�6<7�����z�����mǒ��M��:�ғo�q�X1������q����*�C[�z9Rڒ����ʗ���#x�/9ʒ��
b\H�ң�G\񓩁A�k�[W�d�)RK��@�^��|�(��'|�h�pI]�$Z��e��'K&�ՙFV"�s�g�m.���b�I���%����~�!�[�F���+��$*�T)[�s�I%�''�5��d��`y�S���>;!;�LE�v�sf"N���i�����E,J[�Ej*�>7�\h����}o��}�?�3x_W̛�7��`N_cy���Ɓ����.
9�Pjo��)%b��=��6�HU�\�#�Z���s4$��<���R��(������Iє��M^.&���^���5]�
�k_�Ƴv{�ǟ�T��=��Zc5��}&�E,ȱQ�o<99���g��p������?�7��>e�ʫ��p��Ż������5�cR'8�4wH}�N��7��⻬����Ǉ��_p�լ��ꖪw�Ržj��Q�!iO�D���zӱ"��OQ�|�6|����n�'{ǵ4��[�a�׬BM"I;�c���kRm�Ȋ��"�c�z�=ҿ��?����;�ҷ�.{�Cj���T�qU0�����"�֬��;\<�@UG��ş��>E���/�*�o�&�v=w�@���4
0úMϸ��3�:P��J��סr8��g}��o!5�Mo��mD+˾�bqLq�Uu븵
\9Ƕ�y��{z^<��A+O��[�ʑ��5���
�boy���p�T���^J�A]��Ue#W�p�	�G����:��n�hv�RT8��d;��M�y�( � �Z0�c�+�s���}�=�{�e���Ԓ�kX�	r�]�"(Hn��ȭ?�-�^�K�K��V���d��KT*��o#��E��Ka�@��=��`]p��hBŦj̚�"`z�3Eh�hq�zb�S�G����M)"���cD����E�6�P�DW�D���5�)V�,JՊ���x�|���-gt��*:K�;�y�A{��~�����R���\�J`�<<�����P~7ۑ��G]�k�1?���4�!���u��n�j�$�pI[�����,�W�,��ꔔ2�v��{����Q3E,:�O��0z�L����E��\��
��+cn��Il�t�;{������Ǽ'F��RB4����8i���CV�^�M����ny��C�������8B�~cR��.�1j���O�Ѱf���op_�����d��>c����ɗsǦ�h�G���ԁ�3UH.(�yR��;�����ÿ睿�-�ߺGZop���@�&|��plr4s,��{a�S��=��G���ko!UźnJ����,���~�@s���HY���m�d��z,r�B��T�7�T�Q#Nr�h[�?f��;�D+��+�9�����6?��ٝ�B8�e�۔��u��������n0�J��T������W�x��'�V�F�C��/)�z%������BV$"c _.e�-���BJ�Xf&P�:�T�ȴ��+嚧s�E��Sd��}8�J��`1�D�.ʪ�i��8c�1���)S���1�Q��2�˔��K��j��?�%,L�p������f8�c���Q��)}/jc��L�y۰����!�:��"�WLLs������s����7�|�ӧ����E��}�L�!,�./�c�/f��@���P����[o��+�M#��Į7�b17ǈ�04��7���[~��kK��	��J_c���pn�C]���\UU��u�����r2tVp�q����P����* ��5o}�/����������7�驶W\��|�����/I}J�'־��C�Ф�\Ν�.�4�A����O��mՐo�e����B��(���˩)٫.s�Tb�P׏��'?�տ�4UEUU��O
q�|�N��3�)���w��j�����_�������c�w���Gy���1���	\_=���?㋿��V�e����dN�&��L]� 5�%�K ��t�9�Բ�d�R�e\���x��ǩb7�c���s�AsE	��wH�$��}�Mn�����2���
�I���\����q-��F,6JI81.�3��͑S&c
���\��)��'<)%s�r��	�3����(�"f��)�֚;��'��@���"�[ �jI� Q���ORD�R��хS��t1�4�2�#��	c4ӑM�)f��~���<S�~g��L7�%�,B�qΉ���r<��\�ho0�V'�&$e�]���{с[�t~�5���ʄ.�kzm����ɞ�Y��倞f-���E���r��e����ze���0YNk*u��k�ӖP��σPŻ�ogd^�&w��`c��:T�i�΂��$�`)~hM�{OUR�r��d|U��Vd���}�_�'�=���^��/���=O?��������O�G����G{�.ۮcS�5!��S���g�*ɔP.�$�����cf�ƛ|���MX_��Ɠ
��6�Q���4�L����VL��7	�4(7ǿ�a�Ӑ&��X&����׿�5V��ޠ��~���ﶰ�^����������o�Zo:�Sr؃��2|��_�*&mY��Y� ������qO1��?W�y�~>gK㾱ߪ�"K������W��wi�bY%vM�s�塏粌O���qPz�T��R�̧c^���qɤ*��8)��c�w�����������#��ߧ���s!\�9^��6����N5�pa���$�� U�s���=���"���P E�ܔG)א�������kK�~�^�"0ms�10�,XE/&�gƤ��|N��M����hg�˃=�v�@F�ia�i�IXЄN�Dp@��a�;G�j��$m%+U�4G��+i��������;�9�P�z
�47��ϵ]ߡ����l�V��L���%P�o`1�8o1F�h���
W��R��J���6���_%���|��u���j`����s��K��;�˛���,g�rx�t�^i����� Ql;Ү%�L��k|���{��.��#�2���.����b���	z��`�)s��4-i�v���D&����눩g{ݡ�5�x�.�����t�����Q|ױ}�9���8�%z;�����_6��us;g��;4�s��'�e�g��8�zz>�1���3�K���t.K�s�^���Va}AT;"�"9��njiQ��]?sSL�-O�L��ilȒ�sr�ϯ�A&�1��7O�CSq��M7i��r$�99������
U�v�j7Ӑ�;oSIs���`9ƙ�t���wKL�軣�L�C�	��X����8��s�!"G��t���L�\��X��&��x#M�a����i��e���ک�f�g�A8#z����2jpSЈ���%�!�:��޴��3^W���G���I��tL���4��l����W�Z���7��RV���z$$q����3�?�\�AHj��3��!�����o���ﲕ��yK[u��%�4q���_|����o��]�M�1���A���TU�ŝ�5$P�b�	m
M ��^��)�O�a��©��*8P̬����{L-��:��s�#��l\_?����x��=���[���z~��uLM�-���e�������	�����yYfz2v9���W�X�H��ʗ���T��qK���7/�l-1���ea ���M��(a� �B0Εh���4	�}��׬2	�������������w	��h/8?�؏�,ӕ��sm��gX���&v#�%�l��p.3t�E����K�SS�M�P���a=��$�E�s���p@��D��A�{?ʥS_p��5=`s&�2���BK��q��<���&���m��s�~� 0hf:"�rHm/�c��M�NUQ�ٷݑ�4��I��%��Hb�z,�--"�z��hC�+Z���6օl�Ź,}���n�'��SDS$�ۃ+)F4�s�,Ox�4Y�I�f��/�����ﲿ�#V�Ry�}��M���ez���_�����'{r�ǲgʾB�!�{�]$x���;rL�ۖ���%`��DM�R�XSo�̔A}X�%�Ź�g���|T2+C�kw�*�MmX㕣��?���ѕ��~���T,��9"_���#^N��ϵ�sz�T�'h���ίPU��7��ۇ#@gh�[`�/�_/CӖ��0Is�	�Dh�Mhj��&�iB2͚�����i1۟�s�7��4��o���>��Tܘ�=��R�8R4�>��P����%�HbpŬ85S��Lß���Hc:j#ibF�3�%�������r﹤<^����1�����~�9��6��H��6����,3���9����c��K�Y�~���{`��A�Τ]r�gL�\�!�e�W_78��S�����9���6Zy4���(�na��x8+�3^$���������j��jK)J���,#������������\Ea������������wp��졉��K����R�]J\���mw���sb,�8	�u���JV�v���.��r�}]�aA�2b�H���#d�KB��)O�_�ҤTKJ�$��S�Ū�2�{A;�!/�'�@D�K��5�e����H5ĝpr&���3Z��ɐ�S^��/��3O!��=5�ve¼���9f?���\�l?�ӯ9��P�Ճ�R�ʬZ�}�0��f�#��&�I8�����,���ǽ�����T��p���r����U��d݃z��>���g�y"�[JKԎ.����ՙ��ڴx,�b4"�����GJ��Py�l�-��{oV��*���81�+x@~s��C0CprFc1=&�Z* �66LjF�S�������㶿�j���|X�g��=8W��A�T.���{�Bg�b$������#��c^&<ZH?���TE��8	��)9	�]����zz����tґ����X�-rF4�|��$��JT����{��.�������{�*�$By�Uph�ӵ[R��Պ��1��E-����	<Y�˦«����n˭����a��mW펋�.�78���(����(>wt8*��^S]�qA�}nd�3�G�q��s*'���{�U$'������BNJ�9)u��.r�Wl��׎M��펰Z�Վ�&R]s�vH�qig���Q�kQ�Xi��	*h?}�'��B�fNϷj��hG��&ʎ�|�EϞ}�E����.+����!�S�>8��1��:u��S5[�ꖍV��6.�c﮸��Ⱦ�B�تgU�F=ɷ�%����ӅH����"����Hlwh� ��eZJ�Ԍ?%��+<[��x�}Ɠ���U69*��R𦏤&���kb��#�,7:��h�
�y����oY�۶#Q��gY�	������H%�`Z{�U��'��I����N^��t.<ng�X�d/Q�<b�Z.�[�w 骥WeJpWV��.�$���-+�I�=�z��8o��8'���)�	j���V�(�]�{Ż����nK����1Z�l����*��B38B�HI�. !��S��:[�3���( ��@!�處��`��
��9�"q���hs���:����`Dq�pfr��j���e˨��B���␴���<�or@��	3��5uO�ǋ��T���C%��-X0��!V@���n����/���v��c��/yN����f��cű�\,��y]��O�+_;�dO�]��>E��,���c>|��˧O��ʊ}�,?tx)%h���f��K��y�����	~4b4���M�uM/��IV%+�ǩǫ�/~�<rpoZ)���@" �k����|B��􏪒5��FM}�yYK��j���|EJ��#�i�u��z�R��
V2�Z@��'g�uC
J�$�ӽ�@?^�@P\��FH1ӥhQ�c��cR��bs�mY�j>y��[wo�}�{|�'�{vŝ�-4)1[�;)�C"�85�ISy��������Q5k������K�� �FLsW� �J���Vu��e�E����{lћ��C*�:-¢�5���j��v8�����uU�Ê��-[r�`�!Mo.@w�֘��ZvƸ��ċ,}Sz6�s����y���Y�xZ�:R�A6ԡ��f��@K�4������S~1�i�6̓�r�'ɂ��aO x<Y���f�⋒�H��z<��3�dh��7Z�}~ŝ�6�=����6>8�G�2�(�XϳƱ�`<����a�J|��[.*�+���j5�	��{�'�l~��7����D�(���h2Z��ȩ�9�s&��̵���U�Q�9�pL�:H��&��q@2;h	� ����l`2�����9<��Pc�yV��{nݹO������q��r�r�����|����$��
:��,-���R_U��q��'G�A�/��0�{c���*��(z�"�Nx���<y��^X�C�7��Ϲh8K>�cfd��٪�ŔQ��"&�ȫ5b�BJ��	ΏVDGK�ά(�G\�|�:O��WH��M��g��AUU�W��Rd���=W���?�c��ϐ��<�:�W﬉�~�����	����H�
�x�zE�C�D#t�*!	h�}��e!:e�d�?�]w�hy��67����Wa)^��u \�|���@� p��~�9��#���bG��do�nH�*�.)�xr��(D@$�N��!�(��0
����!K�^Rh���6<���$<y�}? ��!�ba=҅캉�`9D���K4~�v,���%�ąa`�3���R�K������kv�}�yw4����W������ѧ��;�]\2���o8'�ee�j*���ܮ��Ym����5U����)?b��f)H��U����AFJ(�U
�4�Ą�M�Ҹ@�c0���/�D��������vt�:<M    IDAT��0ѨA�R�J3�	-΍��C[�h1&̃�q�oIV�xv�^��ϟ�����Mɦ��]ד/�������6ͽW�D`�\���
K�7�!�}���ĲACh���ȮD[��}f��r��AUm����, *�2�� �,,�l��YW5�>����#*�33��J��1��S�"�(���:��NP1���~M� ��Vo���g )������b�(Q�`�=J��i>k�w	6��Is�>݃'T^��3��
RF��D���$Y��ə��!?�_�g������_c�ګ�������1���ͳ?����^�����0j(��ݖ�
D�))��>s�\�ڌ�64��q���>�я�O��
�8��k@h���!I"I�����PQՍ	�<Z�oLi+�pm�-��$�3����6e�@��~��8�xGw}�:8�XΝ	�������tH��h�W��x��s������;UqR�jë�����U�1�j�Ӷ;C\G��(�V:N)�<l@U��U\�C˓��WCP<�E�,l��|r��!����X�T��Wk..o���_�^H[��-1����DK�����1�1{P����	.g�F��E$W�>��������ּ�^���vk?ƣ)Ƴpr���|{����^��`,��L�� M�DҚJt-sx�M��8���9Xr�6��5Hi9���|�i�ĐQ`Ea���/S�<0>t�a�gU2ٲ��#�j�;���,ȗ5�/]7��#�rl���l���s���.�qօن���/��_�>^p�x��T�i�5�xuE��6�^�ZѦ=�3#I�|�̧� ��V�(j~.��`����d��qD���9���1�aG� -@ҿ:��T�W$G��s��!�1Q_��կ}����A�+|�x���!j���Q���|Ԧ��#��ׄ}�V�7��O���=�3��TUE������ffw�0�T#��_����C6�\��X5�������ן�ʭ;��{�]$;O��T
}�ȕT�}M@�z�7+>x��W��
�_�������{���1��.�	t��p8xAK݂%=���,�c�=��	Xb��K� �5ѧ�TUI�@{� O��-.�ޣ�ܢM����$ M@�!�iZ��Y%�5�L�����a��6;�=sE�&�~�M�9�*��q�|4�+\\d��L��[A���ӱO��qN�=5�3Ӏ���&���y�E,���DJ��!���W57A.��CC�q��s�����g��g����6kT� �R�*�w�Fq}XC��+2#�U�����[�^�Zw�	���ϟ���E��	�0�С|{v�u\EO���1@pF2��j�%J&����S���A�M7��f| u�r��LPǦ���5B�,EC�C�~7? ��|��&�A�9g���R�Y:��K��>=����h����Ao��u҄
4��w�3��;|����'�7��G'}I�4XRh^P[C�n����F/R@fp���U#����9��
}�.�/�I�/�~��U�Tb�{����\I9Pd�I��'��xp�B�	�y�D��� %����0�̃ˠ� �c�G��9�����kw��}��<�}���>e$%�U ������UhU�^��'}���R��_z���/s�wiDhV+4yR$����d����<T��יn���3r墳�t\��\\��]���Z|pd�Fꪁ��^�W;�w���gx"���t>p<ן~@��hL��Q�yn*�.E�XƳd���d��:��*��$�Q�-3����9#|�O��4��}�����2Y蔎~�ȟ��������b��"/e#��^�
j��K4�e�lßK���=F��T�?�i�.�!�b���Qt�k��g��S }=?��<
Z3���X���,-4mw�P���b9K�}ܲ�wH��lV���$��xWXY������Į�,W�m�651G��s��zRn�b�Za��Q��!��ދ`��S��8���td�zB����/L~z͒V���n2S/],������e}��ִl-�
��O���a��d9k�d��9B��62��:���g�g������j�፯}�6�.�<z����^�|�fz-�˖
e��m��8�}���CD�W~�k���׉��%�	V�������'䂌���O�G�Р���<�*�T�'d�Z���da�����k>���>@|����P�LG���5��yU��2��q��������9UThV��o�֗D�H"�P
��/� &�X1�I�O��k֫�\'���6���gU;���츾�Y0��O=��:@���Z�+��p��l�Q�����UR�D	�q�{�P���
~��c����T�2sgR%b�[��b��oے�bܚ��k7�B��YuV�X-ۮ'�[���!��G�tI��7ͭ�Kgd�|@k;(@:2
!q��+tv^���~<7��kD�*�Mx&�;�>)5�-�b(*5o��<�<�?�K4�E��8�x֡*�$o��(�Ij��cN��ں��CE��^U�u �$�/���kѱ�z��U�\S�*�uv��ytM�d�Ư��/��t~\�t
 g���R|t]in�yMs<5�G�NM�c��4��C���Rg�5Gܛ>c��,�������M��#��ك]�9���ڋƼx�p���WOS�8x��Ѫ�O		���$8-�y���q���O�e�����Q�������o����7�ФT8����o�uR�;�ŏ)4� �/��gR�r�]Lt)�EX�)a���	q3 ?v����ȳ�>!^=1wAU�>X|UQW)EL=rG/#�%��=����C��G�E��Ľ/��嫯���z�eߵ��̫����'��~e��D{�N�]���œrO��S��~��Kͭ�%V��Kf�^[Id�H��o��������|�w�C�Zq��<�����^�Nh���e�)�IbA��A�Z��8a��9�����\𖡠�T>�Рs�o�%�Dլ�u���#>������s�H����Y���+b�ߍ������.�)m<�z��$�,�9�@��i~M.{�Ua,#cg��7T�^*�������ئ�/��<k�L���x�r��u���g�Zz�E��Ex0��v� ^΂��t�If@�5�O5�l��Z�WHv�{;��&�?�NL�.Ym�ܠpM�>~�>r�%�b�=� ���!�$)��oQ+څ3�9��>+*_C_o
Ꜩ�V�J��
�OhT#�j��":���P���L�BB6�ɸ�w=�l�}P|vT��r�Z�L�۔XgG�+�ޡ�W���-����~	�����%Bu$D	\����o���,R AR��5�҇庒�~}Q�=�?���X�RG�J��&@�l�5&3��CD����� �L���5Z�i�P���Zko�K}�T�Y���;\G���?�:%��oj�EX��&�ڎ�w�Α���\%$�C�����#Ǟ��^3MӰ�n����D�.y�W�&��5�k�I�H�=�+D* �z�fֻ�*��.�\Wt�w�u�xR��=�y&���U�'{vx�������2�����,�>����W��<��U#��9�����_�����a�.�����
�ЧD�B�#]�*=�Hū�ˆk���i�h{��hE�ޣ��Np�.� ��<EG-��H�g�6�$�#��m❯�����7���x�?�3����ZwAV���O-=~A�@ސ�=�ۓCǣnŽ����_�u>�s�����C����c�6�����=��
�I��O�J���;v�ҭ6�*s�:�O��~�C�;-W��ʯQ��iG̲x�hh����%�(}��Q~��1�o#���'�Zc��q���p=Ƣ,�9s�B#�/�l��1�܋�*�
%%�X�Zisg�"��r�adFK��ar$=XJs]P�N6=�'��9��m��Мs�%�Hto���z@�qNY�}E﷤�� ����'\����d{0�`�!�UL�ԳA�q�8��R��"�YLHN��
��<	�Lƕ��s|�u�ۖ�4�D�z��t�؁�I��7����-�����|gC����3?��>@�ؓ�	��6��1�7�tc�wF�6ka�m���Z���aS���o~�M�z,�5�R~9�X����,<�Gv)�KV�q�z�}KK�p�n�����M�/Y$�������|��MS�R"��*��'�6MU4�i�|M�,�������P���<f����g�o���֪�س�z��9MmY�ǌ�Ү4�*x�������*_~�m�Wy��Yf����"8�זZ*2��[�ܾK��k<M=�S¦Ƌ�����l�9<��泋iON{������'��?�Cx��~U��o���x<���i����\	�g�cs��l��Y�D_;��q}Es�z�_�o}��zܓ��|L}M�Dl;\+����d+X�DE������/����=��O~J��)uj�ԡ��Ǽ��9<�����d1u]�$�.Eb�E^%�Bz��N�I�+4�K���TT��d,�d�`�i���w8h����M��6��9��YKG��p2��&H�mF_��G��CߦBҔ�h�=q1��r��U �L�w��I7���Ƴ��c?�&�r��g=9���� ��ob��/��)����<��]���~)O���4�ab�~�'�KI�p�QJԧL��L[�������e�T�(j�<@��ggi����py������ ����|�K~��"���y��T���U>����3�UM�+nݺͼ ����c���L`>��χ�M�Z�����|��g�\NTάZ _�q��hm��p熠�L �>��~�q�o�U��X��v�����Ԥ8��%8����d���1�?y��xǭ׾���o��;��h��}˥ `u��h�#kO�\�;\����q�B�ʭw��W���K|���ʪa��+1SB:7]��["������#���w�����_�y�u|~̣�����Zi*T��`��-���*W[a�U�r���Dý/��S'TW����Az���B��J;�� �s���Ugs������WH��YY���� �d� H�y��J�LL!k�6ׄ;��\�Gh�)�q�Q;���r����2�y����v�wA|���M�-�lu�䚥{Y?��]����������	�$A�۸�4}On�%�Cȉ��'��9���93Ec
�;�i\Kg�t�
Sw 2���������H�A@ 7��qB�&�֦Lf�q�Es�8q)��Db4�����fS�@F�RJ8�R
o����ʱ�9N��M-
�z�!0G�ZZ��{�q7�*R���"����^���B�b�{N}���{����t펐O|�Ï?4�puC�Z j~�A�6���7��5�˹�>'���	Iw�b�ۢ�*�ۗr��G�.3N�������i�'��sڇO�l.���6�2;��w�!�Г���׃����|�'�g|�6+���_���:*�
�hƹpt?u��H���������Ct�������?��g[�X��o�._���.\���6�.�X�N�L�p>t��@t�ٱ{����@�p�wy�o�����&��>�������!!+�Ԃ&jY�}��>�յ}G�H�kv��.qs�_7���\6"��ǚs>c18�����	��R̈a|Ľ�C<�����}k
�,�i�b)��V\���o� ����{�ݎ��9���m��ڋ �8�ʆ��x��(�S�4
r"d�L�2��~/�ї�O�Xrڪ����3�r]�x�D���!��%\��Ǐ���b�Ss��5��9=2�����l?Lg�鈎�4�C;0�c~�~���_�}�tN-�~ДG�����sL؇N���;�'�5Gւ	c�;P�j� ��A����P�"9nK�4c�=�W�"��@%&I�y�˼�λt�@y�L�����ub6<~�9z������{_[)ݾ��D�k��tY�F~~oU%�LNʀŞ���,�>߀`+���aÏB!�9��HrЊ�[o��%1g<B�E�^C�9,dӖ3�"�*G ��?��_|�������9� �؏ź�k�4O&{4f�>�*G�Z���Gtۇ��%����5���T\i>�W��jV�5�jE]5�}�Ʊ�o���K����7�����C��;��Ϣ��y����'G"�'1�{�����Z
�[w�?��~�;���k^��[����O�>�U��#�<�7Y} �:��`��~�V6�y��֌Ӗt�����7j�jn3F���,�Xa2 t	�jE������ݖ[�`q����P[�/����eO�%���ݯ|���|��پ��Wb�!&\���x��QI�=g����~.���jY(�P��|Z��f�㆛�O!����~�6�O���p���5��司��3�i�F?��0̳ϚTs�A�d�΍��S%p��vt�F>�k�(�t��HǱU�U�!g`������b�g�|�	:"\��rn4����5��ξ��% �O���u�j�2�=�?�z����68�p
"1gt}lqU Q�ݎz�fǱz�>�� g!-ޣ/��6��M17	/����>�﫦���.W���2�s�9���Yn2�O��&��jnȨO$pa���������<�6o}��������zb~��C��V���mA��9QE��I��N�G]��>�r��(�G��~���mۢ^�\�\t�U���S��m^��/�6���;�8�Pr^g9M�Ѯ3��n�������Bp���<���v���;��?������)�:���y�KZ��Ͼ �m_+���c���7~�/�������㚧������{�1��v�Ka�����͵�.�(=��}/��o�����y���'�}�z�s�k[�(�����v�n$�ȯ�=>A���Ɨ�ү�M���h��WO�R? ���V���\�^��.�\e��W���o��k>�����Xoj+BT�!�	���D��t��rdݜ�с]��TS��Q���d .��ꛄ��>/��-���!ܰ������{���O��?�駟�i@ԡ�,��s��ߓ�EJ�[q�O����ð��#�	�PAϠ4�4�s���X{�fI����w�̬���4 ��6Vn �EC���LI�-�'B�_���3̄�Bc�c"<�4�(�(�$n"���h��ܾ[U�r�8�YYYY����ڲ2O��ٟ���s��\�i!em�n�6�%k&�	<�R�rPT�<�H�J�|_��������Q�����_�~���;���cu�s���,�Wl�(%(�)�P�����Z���[H����q7	�?��[\��y��g�N�ɋ�
A��+���a����nֈn����!F�:�Åȼ�����E��������S癆�W��W>:�A�zTL5�A�J8�`9�bFF�g?���r�A+�N��s k_m$2A�����AU����vnc���~q�,����e��g�M���4JǸ� ���o�V�ݟ���?an|BY�L�z�/��M��}���]5�֒�"��;}�omW��q�i^�����}
��c.��ſ����&c)�F!�(M�!�5��h�ٻ�W��(H�!�}��l<�f�0��}.���H�LTR3ɚ�w�լvg1VR:Cr�Y�<�z�QŌ�+�����	�Aym�VG�-Arɉ�Ԡܜ�ﾆ��%It�
����c�B9���u�uL�+����Z)�$|eqe����Z��~�^�h�R ��g}j�7)|1$ַ�H/ڤ#	EAug_� D��5>�ƽ��F(�������c�FX��j�}����K#�/��Pk�p]**�u�=��MU����dF�J�ެ�j�.�6J�Z�(�ֿ+���J)<��*�E����Z�{�?�b2�B/Mp��j�5}�:��9�I��bz���;��J�$JG)�uJ���M��Y���&vq�Z�`Õ�    IDAT@2�LZ�a�g�}�y�ls������kw�����I�>�k�;j-5�)��yy�2���7�:er���9]���8�}S�{-����
�-؂�?`��mB�����:�����i|�r���Q��=�JIt�1�8����^���%'�~����iF�BT���8_PUs�L��m��%�c����w���?y�� f�����SO��|p=�<Cs�nn��ٔ3����� �dLu�}~���Ov~���L+�2����lJ�%,�)�ir��Qy��:F�������|�m�YŶ�jD9OaBX�z�{�d�P�@������,���Mv�]��s�R�֪��Z���X�_S�>���Fd)NBb�p�T��*1J��!2�Z����������<$���j��T�r�$�*�Q˕��ߋv� ~=s�WEH�~�c�}Ai
o�ޓOV�9��u��7}�q��J�R���u�a5�X�nU8��b�:�G���F�RJ�JP��-Q��e}ԋ���;_Ea2��bU��"@�ã2M)J�j�LE��	FEk+,R�-�oI�D�ZEbe��}��m��uu���t��m�<ʃt�+bQ'YD�'�)2Pلl$1�!�F��u.����M�ed6IU����&�9�1�#X�w��#XK�Əc���D�K=)M d��)���H�	�n�Zε0cE��c�g�(F�&$�"qX�p�0�<�����.������`�z "eB,s*��EK���F���p�kq�$�F�n*�5�흊0���� N;f̑#A��o�g0*E�ĉF@�,N��č�)b����@��vR<7�I�l�1���0�u�<q?�}�-+�*����@$����mM�Ԅ<�#���B	(5��ܘ�\����Gd���^�:�'�Z��i����8U�]�,q��R'*ly����4��!������{I9Ҥ�\��ϻ�������k���䗮P�Y�D�"�B��r5"a���pY��*b�{J	��!�.�{�f��=w��?0��+X���4�s��I�鄢�Pׂh������g���g%����rx�,g��,�l���0�rl:Co*��)F@ad�|�v��I,�%�Ra�B�1�,�$da�4p�_2��˨���U��U�U�2̣�,ηM��9���l	�b��0uY2b�T{�T�&G ��S�1Z��-�L�� j��uLU����*3�Ay�I#`7�saۧ���s��)Ey���D%�2�]� u�ͺ�J�\ˤ����)D���>�w/BE�D��S8��pZ3�6H�&y�蠑>�!��R)��xvu�5 k� !��� ��!�AFDH���*�'��@�E dߒ�ڽ"H���(�̨�2�0B��$�� T����E,D]�k@��x�s�q���S�f�FS��	h���6��d]_��	�X�Kf��J��������oYYdbVҿ�` G��e��Q��N_�m�G��`:�!����e^��	���Q�lE�k_t����Ǯ�0tָb���`�̴2�����=O���O�p�DiL")3C�(D��,p�р]Y!T2x������v����he�_�A�JP�<�7w�Z�T%�s�%����	��}�}��6��WZf������'W��

/9���4:8��[��2��Q����jF�V%R�i.����������S_���#߻���f9FT����{���$!D��t8B ͣ��	]����gs&�3Έ���)A|�5�n���66E�����7����/�"�����:�g���1����5C�xDP5�YmMp6��[��ן�o}��܍O���/�Zrn����121��m¼�z�͎���'��
��A���tc��=�@}���ɄYp^Q�=ގ�唲�Q�C˶� [���E�4��՘�<ʉ��a��]��=�!e�5ro���\��ۼ�z��:�~i�E����:��:ȭI�t��ꃥ������wRJ\��@ �k!JEs�V?��h���������D��V
�d�����%k����"kh�2��9�? Cl.=d�ۢ��n��⺂�-�Y��JK�j��Z��yԍ��k&�����LK���Z�c��-�>zk����
_%�c��Dw�����kS
�� Z�s4כ͇�h������*JTYpp�r��9٦���Zm]�X�T��G��Qf��D�jl����#�T�Q�*�lʠ�'����|���g�E�a�#�]&���ИmewgQTTA�y���E�D��1�	p�.�/]|dJJ)���Bx�������՟�)jr?'^�:a�׋9c��B�Ob���
ӫ+ߝ��ϥ��"�$۾��|������Ԩ�u�ch/u�rfl��T���>��w�v�%V���C�i�:�QTH,BƠ��*G���=Ʊ�����U���7������:�A��<��r%���>����Bh6�>͹/}�
�μ���Co��{���x�ŮQ%cF�fb�l�%Bt���ªן��ա�|�6t�\��O<�����wns�ױ����S�����.�o�;4�G�k�X�mB�$�Z����ֶ�����(%�ֵ�4V�~�kI�y��%V�n~���>��q]�"������5�(Գ��ʄC4@v3�h�,���z7�.ш�4���EbJ�#�Ng��A�bw�@�k��\g���'�ߧ���"�#QF�|��%I��檘�f���Xh��
���¥��8�]��hj_�����P��%| !�*�_y�>��w6Z#�1>D�T���<޹�t�W�eh����mCX37��ֵ�P/w��.��SlqȜ�ѹ�8��yG	�Dw�uNjo\�)w�u.�0���Gos���x���<�ŗ(��2��I���>G#-�L�昮(?x�)3ax��������mL1݌�|>�V� �JǬ*	ac!���ڒ���B�Q�2��F�^r���I_��5s��U�RUX�g�\9�]�D#�ܲ���u)c�\/9H�(1̽���/rߋ��4�M7���ט^���B�W��0�	1`�>$!"!ʔ�O|�cϜG��n�n݊.��ؒ@X��w���2�����29u�9���޺��CM����G����Qܺc�A����ݼ������i
��SЧw���ں�����:�7~"H�o�$�)�.�T��&�v�9vt�P��!�ꀸ �@�Ȥ���}~! q]��ǁ�+!���}[�O_���ˮ����f����ҹ!k�N5~��_��x�#���iJ�y����y�"Sݖ5��g@R�N|嫘�m25�Ō4x��T�cn*��%�F_��>�n�"=)�Epc+}�G����}��јE�C@'
�w>����!I4�+�S�u���%;���֭�#��!�͘7��{-�ad"��a����ipxeH����1�|��4����owLʋ`�-�3������ޯI�'5Ǐ��DG���l�N��1?=Ib-��mnq����0'�5������䈇��M�#O2�:��N��1�&#0
'$��0�F�ٞ+F9l�	��(�
�(+�XO��klHp�� ����ȲB:Ɇ<Ɩ>��e-���Z�W�G��-@u�4B�ʔ[6�{��O<�Xyn�����ۧOGK@X\��X�d-\+��ף Q�Bu���{7���s��7���l�u̦?F��z{¼(9LF|������=N~�2�}���;��:־rV���1���?����V=��jUU��$Z!L��{��:&߯���.�ِ �d)��v|��JE��j�Q�|���f���o�9���C�":j<�L9~�ľ��$I�Ib`hON_���QLe�C�21]��!��k(iV��M ԝ��ؽs	��h��h4��ߝ��>��u7��j=Si��a���ٳ�<w�Ys鱱��QSn�|DL���e4��_����@k��KV.�|H���x�'T�`ZQ9��M�Y)�	A��CsޞS'nIa[�O{4�55cb��F�ׯp��/�v�Id�d|��R�X�}X];�y.�a9��{�x� ��k�1Ĺ����ؗu��n�\���yQ M��&u��sk�B*���	7~�3&�.�[6{�s_�=���`d�$MЩ$d*Vg�-�����NJ�D�dAc�����§����6�u߲���,D`(mb���KU"��к�L���Gj�L��p�Ԅ�� y�	
;c��K?�;�+�Ʌ���>�H�ø�H\�_U��*��!�x��g�2S��7_��P����AS�A��R�M��ǣ�ۏ>�i����?D9X;c�-8Y�pM8r�U�ٺ�ۖ�o��� �6��GD�~=y�Z�h�CM�:0�֛��h6*
�!���(.�Z�=9�CB�����������-Ʊy� �o�w�9��4M#���5vͰ��e���i��vd�D��K�	}������C��P�ʡl@�U�\K�E�4�C}Z�ai|����Z�R��V�F)���{!8������?�MRD�����ۜ�r�Կ�u�`����j���.*џ��7��:H��C�@U�TJm���'�i�}:�cլ���c10~w[C����������.x�pl�S�k7��2��!�P����0?`�-�ܣk���xf�2�,�������Y���'8�T['�u0N�ye�k��XFU�	&KJ��@q�d�`l���1�_�>���
�~�l��[���l���9�,w�c�Z�Ts��L3O���U��(Cld8�r5?�%�Mc��Qw���T'щ�4��$�L��^�a���΅�Hm>�l|%$ӓ��ķ�[x�sd圛��1�o��S�b8.g���Ѫ��m��*=��/~���}���Q\��h���?'H�r#z�q�J
�#�1�a:�oڴ߾��mC���?M�����C e,�H�����3�~���C4xM�^{��u���uiQ3���W���x�&������!�g���t���s���bY�S�|���
�����}���E=�{i}�a1 ��hC�>�&!B�*���$HRc��n��,[�1v	��d3�؇��Oj�fB`:�����;;��ὧ���[�)rlmm��F���3��ώ���X�kZ���1�7X��t�ݢ�4���#e�J�����T�et�꽬�.�<0`�Z�F:7�;�!��wP�	ac��?ǹ�z�b-:��1�r�Ս��� ��mQ^���/���g���SOs�N�i��*Te�$�� ��r��*�:I�b�!�ۛ�勼�w���k0/�N?�3��&�gqZ������I�1Sɶ�TCT��i CbrGR	DU�ʂ����>bں�����UxB9é9!-�XL	�Rk�V{�Z���K�� b����g<���a��W����������Q����8��e�*���s���0�68��9�q�����]�@�u�����J�DEYM��%,����Pz�1G	۟���#F`�
����1���{0^�/Cty]?���K�T��O2�D�=5m���Z*[��r�1�n��w+Zz� �Q8b����:N,c��e�t��V�mqf��Wߥ�}�n�j�"u�}�du���`��m�h��}8�k�Z��#CL7S5��d�!�)N	lph���^ͱ\PhB�CG-埋5�j���:��{O��`y�&`�	{���R��E؜���+����������|��WX���<���O�S�%H�� (:���7�!@P�ܻ�I! �%�!e�)���l����Þz�2/�2�TT�t�*�idI�`h�N��D�k�T���:�)XWC���K�B�uUk]l����D����]�vq������l����ܿ�JS��L|� )�`]I)�x�
)TG��A,,����S?%57��6F(R�=�4�3Rlh�(c4� �$��<%3%�9.ߧ:�%�hW��gqe���I�4�lm�P�_����o���T�8�����d�s�l��W��p&��,G�RD��(-�8p%�5/p�C�[�&�z��Ǘ��F���jP���)8]�A�>q�RX�
X��A�*�p�P-�s�h��2� c����}o0^�a=2��.K����/�>b�`����9�ׯ2+��2�y,VTy�T�c�ؙ��Q��
4c��XH�-=|�o8��s��|��ox4������h/A�t;�A�0�B�zM��H�`��g��ǎ������աŸa�1Ŋ��jه<$����ܫ6��k� x�(����P�8���&�x���&�$Gp�P8y�y�q���f²u5�U�v>�����{���m�`%d�O� h-�dX@i�'	�L�L@�=�<�L>�؜P1C���b��R4>�D"}�w_���-F�ŴZ�[��%RTH��b��"�J_ã��+\z�J�Dh�4qO�Z��%��H��FF�WB,�eE��9o!�APZ�ts|b���� c����5m�	��[��i��v�B��U�W�����nnQ���^��G?�{���ѦqO�$�ٖ"@>/�ۻC��̕��$F�\D�`�WQ��cڗ���C�ꫦ�e��O�2�v$����ػy����N�G�R|L���AjEс�m��O��GW�鷾�b�����߸͛?�)��)�C;��cfJ�pH �Ht�:Ru|�+������Ûש._���>�(O��e�*Ì��ST@��j�*��j��E?��(i��dQ@0��Z�t�������}{�2��&�}�T>�ua��M��1V��DL�z�{u�����
��b� ?	�%߭u���]5[.�����d�:���"��Da�do?��{�s/�.ũ�I������x�T(6'�0h\Y��_��s��iM�N#xZ[r�6�?M1�PɊ��磋o3>���ٴ�V�7d��?g�JI��:}_���g��6W.����G��I��ߣL�G=����.�i���D���Rd�)�q��c��ӘrF��G��S�-�¡䪵rh�������V��V�
��(�����<���8��9��;{�����U! �����+������[W���?,|��R�~k���:��Ki�g՗Бhd���y������;f�OCSUCк����վ�ja���.I�=���,�ܕ�x���h�1`c�0�
qX��� ��8W E�a>i+��E�R�� # zeȠ����M�l�D Ձ[�����ER��Z�,w��c3"�����@���̾o���}R�L��s�yZ�*��{��L��bs�����)G�Nz�X2��8_2�Z�>�*����`9��c.��)vac���}	9y���R�
�Ā%�h3Ai�v�5�fr�ƒ��W�H&����s�kQa�x�1>��?C>��wgdڰa2�k���~ ���6֏q�i�cnY�`i�7���r�߇̂C���k2�bns�PrX����2>�<O����c��G̒�\��?�r]y��*�/軛���E���t�����(fE�?�_����� g�L?~���%��`Q�}�34�!K�E@TJ�l���O�*��+̯Ȇ�UF�i�ӽ0�n�V���+����ғ{˾+�㔓_�<�S۔W?��/Av��Z��:����}�?=�Ueb���[���A�����m8��L�����p��@��bj�|*�[�s�g��}��(�z�~!Ze��6������V����S(�6n��74���<�F�Z&��İ���� �F�Ie�^�+Q7APem��6��*x���4`*Z����\>�:�e��'�x�� G)C0
�.�L��=�̽��o@=�C����H���t6�� )��D�t{�
�z|2��ڤH
O[1���C�5}��?4�G���'t���bk�rJ	�b�2����<�;@n.�ҭB����{���=�1�S�s$�dÕ���I�=n�9������^b� U�ʗ�4�*
�l�b��~v�a�D	�R̦H%�J��G\��������ȗ�Σ��o�����AIK}U�    IDAT���TSUC�6Bd�1�VՂ���
����?]�ߝ���)-S�� V�O_�Yg�Y���Z"�~�P�)��ٌ���y���������[|��̵_�L&ʘ^Ti��~�^�>FK�mB᪂Dk�6TƐ�=Ov���|�7����3RLt+v�6aY�ij�Ct���u�d��p'�p��Y9%�%
A2H��Y���wi�%.�ڏ<O	�)]��m��=�������6�ˈ+���}���}m�z��w{�������J��3l2f��}�Np�ݷ��˟QJ`%1'���c�?���EkW,�;��F:,[S��������Ww�V斈�E� �n�bOՒ5`��'�C��Q&�%&$:�L-G�]�5���|s�ƍ��k���ۚ����3�5�uz뚖��N�U�jM[9�k��������3�1;�9�*�P�{���g���& gi�:|��Et�څxR�B�] ���%�z��B��D8��?�ݾM��y�_~�����;�$���!�b�(J�"2���b�����l���
�{�����~�C�x���>O�}�	��Nbk]�D��4�y@�$�`���z���_�ٔt��}�Kd�=@1��y|�ƣD`[�:�E.��=�U4��CT3*��ȹ����O{�(��������`��qn�i~8���e�B(���!h�W�w�~-�K�sw�e'�pu^��ݫ0�c@� >{d�1�<��z���߳��/����E���r��G�d�ǔxL��>V���
J[���r��:a���/}=�z�w�n����a6]��F[b�+
I3��g_��#<�������s㢏6�wwޭ2��o�k�s�3���T��Df�̘Q��XN�%p0e� '@ؿ����KE���#�y�o�~�uTg���F�z&�<;RP��1

�	�d4��$���'��%s�)k���}�h˥f�����/�2허��g��e!�%(�����|�޷Qj!?��G�`��{�浟>��}B������ ��'I���VW�Z'��Z�]���*���Rz,�"gS�?z�G�{�o���������#��bV2����ݼn���Ll��c��ƆK/J	F*���2Qq�7���{Xk9��3l>��� D���������F���n4�����_!5i���n��/_F\���,y�q�g�d���t��>��{ѱH�J�[gK��+r7�����l?�4���7��LmșMw��y���L�yw�0H�P�E"�FAPy��ƈ��x�Ʌ����/��>ˉ�����;��N�k�m�1�������)	^BPD�`�)Lgl���IJ�kaq�
���%$��p͜䁯~����O�:�dv��W�{���M�~���-����_E\�N�D[��'t�$K�u%̊,�T��A=���6:����K��̶��} ���Z���V�'I�<�O}��_z���o�΍7�"�����
=�4L~�����t[�k$�V�J0s��JAB�T�1ز�9:�n}���{�_�9�1+E�p_����#c��B	I���~K�b/8������ۿ�/V��XT��}��A��ի�P�P��hj<  x�
��6�,-����m�xibsij�u�?)�A�Y?he��D�J�RK��L�2�$M[D�~�m�!��^6�
*FC����a����W��W9{�a��y����L�$�b��0
]kd}M�}�R[�_���bX���%:��)�'����KLo\EK�F�H�fd2���ɹ���,3�~���p���{��<�%F(DpL65���w�g���O�����<ơ+�d�u����z��H�]�H34�)H'���~ÝW~�{�Y��/~���8L�!�b�I�)���4��s%�_^*�WTsG�-��|�����?��v9>ɳ�ξ���l-IB�CxDW�� 25G���D}�P@�:⺘�|3,��e(C�!�J��q�����w������5f?�>���?Q�y�LW����#28,�X�^�=�1):1�Reb-��Az�3<���!1��m.��{\���Y���üd��!��5߇�D"nC��1g�cc�r�����[o�U�H��xi4D>�[w~�)6��{})%��d&���z|���4��'Q�#�5"�S�+�\e�_���Z������\���ڸ���'	b����RB��9���<���/}�{eu�7
�Z��%~)Œ�ѿ�P�`��(�����~�e�e��3k���+�����_���ύ��B��7χ�jzQ��jR?��;X넖��G���,e�f([����s�R�J��ױ|�~�.�h5��u���v�W�Ǻ��0m-���Β�9�CY!��H%lLRaHQ�*�l,j#d]ӹ7�]-��ߡ�C�~H+�?[M��b�xd�}>|�g\��I�~�s���)��'�HRm�� }�f�cRH��t1�\MО����~���u*�0g���^�m���Ul	Arg ��l �z�
�(�c�Glʌ�r�D��8A�������z���1&����^ ��b|d����4-)Bx���8V�cW3����4s��v]ʅ��n�(!"�@y'�>�g��?E�����Mn��*���_�����l3Õ�����y5<��\w��yIU�Q��i2y�<�¿`ی��_����9�>,�6ی0�i�"D,1��&0�g-
P���ڂ�U��o^aTY�G��p6v?M����3���;�#Ӧ����lt������SOn����V��I�R�R�+kk�?J���|ͯ��R�2�1eR�#�������"}L�N-�u7h�������"ĂO������=cFR��f��ī� 2���r���s���h�*!�D]eQA�h������t�;��t�N��&���@�^�+�JP���b��h��@h�f,��j-��8 .ԩ�%�H���H�b�:֌M����T��IB�M&��f?�E�=��Уm���;�(�LB���6�7��hU��t%bs!�m�v�A���_�N�Eᜣ,s�P(*���Ʉ|Z���=��/sd����C���"`�g�rB¢��$�#"C߷R��j���:���TY�M��P�I�䁛���*\G�Mr�qmU����p
��� �G�@"%Z���M@��C|�XXR�(����C��>�?�s�W?!x�s����8�3��ݨ(���j����TJ����ڜ橰��ȠI-T�)9HIr��s�q�ɥ�������>���yq�B#u��uߺɛĴ::���y�R"�CHK������J�ҁ"xE��.�B�e�T��]�Y�rѫk�Y,��~m)%F)R	���o��H]c�տ���/~�d#��fL���ɂ���(*_�{�m
f����k��eC�������G?O��qB6e��W���:s��o�sLl`6j��B;&Rj��Q�(A�#���f�D���=�8�[��G���3����`��-aAh��56�B�b���a�� ��E��U#��%x����_�V�)f$ڐU��θ4��=� ���a'#��p��O(�&�	��"�$��m���u���׷��$.�g�2E�|s�=��y\w	hc�����)v��7��z¸4LJ�\͙�Qe��>�4��"4���ԡ���`آs��Z��x�Z(t\@8Oa�/�* \�w"xJWR�X��y�@G��H]kAj��(�X �񷄈7��uI4�!@�qߺ��.��	(,a��P��w|X����B;��J6����C(j�Bgb#3�%Ҙ����CS绵&���5�G�}���Y06<U>g�c����ǏQ\����K�V3��7Z۽�y���f����<�J�>n-��_�5���y���g_z	^�����aT��9<`4�%���Z�Qs���u2Yu�S��Q12
� M��r����i�Z��o�!��6���3�7�4eVd5�uSl���| 1��5Bj򼠨r��9�����q���m�x䛿ǛW�az���N��I� 8\�p5$�ЦN�0m)����]��$�³������]t6B޾ƉNDw�֭�n;ʚ�tN�A-�w��[ۆ�x����W.q�?�g�?�%;����
�-ib��K^�:a��B�(�s�9���5����T�>��o2߿�81T�$/k���>O���V)�+��F���u��>��3��j��_}���PB�CI:Qv�����{}���[�k�w3(CmQ -Z'TeAi����l1>y?�gNSPp��9�t�1�$ep���9�2ѵ�.����~qN�o�|�_�O/�L�� �砰����?���J��=2��@L���#�v�TA�
!!�\�Bͬ# ��\t�%Bk�i��r��=◪�����U�!v���ٓ�{.�˲e���5��;��pr� �!h����ӗ2[ԡZ���Bn�� b�
вK�	t�+�ןWM+fʥ�;�M0t-W��M�s!#:����������������F2�r��LX�R����M2���Ee��%����Tv>����E���O�羧���c3�	Af���������u�gVΑ�b�������q�����~�}g��/���i�b3���ǚ�5�d���$ea��DA�+��1���+�����=�͔�_������~�#�C	���#@F댳�y�CcR�s�XT�٪�l||��ۘ��d���4XS],g��-,�w�����w!��۪�8�O��_��n��{�{O�w9��Ϲ�Wߥz�uF�)F\Y�0�~�q�?�E���</I�B��r|��/~�G����z�vz���Ӌo��9�Xk�mA�*l5_;-�ESV!@U���܎�'��BS$�\���o�D�XXʢ������>}��C�7L~�r�4�#�T3�X$U.P*Qw�\���adZC%"�F���~���n��n��Ex�N��B0�s�I��W����_e��%��@�X	�a����}��)��{��>�5>}�EHm���ǂo�85�oz�.�FI�
�R��d����m޷7�h��9��8km���
,��	m@��=�_�ڐ�3�Ѻ��� 1�JxT��w�৯`gS\���3�!G����e���]��J�B��QBHZX�nU��l��aQPD,�d��b9�,XǴ(�'#|�[��l�ʒ�U|�ƾ���6�Q����1u�8�jN�3�ͧL���M��m��ϰ�d���'����o֨�`�FML��gF"p�hn��\���M+��)���?��K��U[������Z��D�zc��ؑuB��&ZJ
_�vLƞѦ���Nb������pNj�|K{U(����`>��Qs��O�0z�IM���d�����rK}�P޴hޕ�
(���*�l�4��FO>�-����y�o�q���عC��f)Ȓ���v�imaN�'Q� ���<�l>�w����l*��1T)���7�Ǩ{���6�bM[;�}fL�$ �3P�9�b��8��ϦQx�G!VE�x�S�����������ޭ9	�*���!;{���J��7�·H�%��� 8!b�w����Ź�%[`]��h��~)]z��Vp�H��hQ#m����w_�抍�ca�g��θ
@�i�1&j�,����{�!&߾jM�.�BH"�����Fб �A_ vDI�vroA�4ţ&���'��d���ɹ��o��\����&�q��$X<F*B�����b����T������C���(����H��9�HQ1߹ʦ8+����o��p��lBB�0��{�>3�o�!"�����`��@e%E�,/��Ƈ�r��&#�����:�<���Zz�t�ԯ ��C��H�ɒt��X�,H̯]����}��:��ϱ���''�!�y�c9Yk�RM�u[��y���GVi���s�
����Eyա1^�u/�g#/��E[�F?-v�КX&zk�� A9�vT몂�/�ms�@m6v,���#�H�6�sXJ�W��3�9���H�(o\��/~��|�M!�	�g�h��ከ���ue��m*8*�ܞ��U#N?�[g�1��>~����'Q:�0Ⱥ&��������뎣�a��R���"���
�z�)>��/`6�|�b�Kb$�{*�Q�/ӟ�u��g����Z \��9�3�5!�\�W\���k����Rd�+����!<���Z����ߋƜ��E\�t�w/"_[d���Į�yB��%��� �0(4��]�������|�����.M�zFލ��7q��Z_�w�=^������UL1֑Ȅ��3W�J�� B�:�,�2A��!����{n��e��{�����[�����d�p�/q��/q4R+�,��Y�:P�;fw[D�g\7�]�;�D�V�M2l�qʭ�?d�֫�����O����M~�U�єX��fe�c�SY�b�O�pEI �"xA�W��3f��������.��<���y����7�ȃ��F7Y#QA���P��Wy$	R
��S��;mW�^J;0�vtj]�=Џ">j�?��?_��>im�#��<��<:���J�J��m�gj����A��M��_��o~����=�G�r��0	�2/(*�.�P`���{x�� ��1qKJ�g0�O�B�\���B3���Q�%epH���G��:�%J�%ũ��%�a��[;�i��"%�М���z�9�
f���������4�hi�52�U���݋�Н�s)���G�Ί�Ҟ���7���>yTUｹ1��5��	 @� 	R�H���E�j#��`��9���6k�7dQwyI�	�$� ��`f0ǻ���<�CVUgUW�P�/*�_u������0$�R��$U��R�e(���z��P��*<M���}\����mr�Qi�L�~�7��I/�O���<_	�qTY�������}N�5$���E��ĭ ���Վ!e��Z��
)WN^�2�������A%��q�խO��0��w�(��:��$�CX�-a�u�c��B>P�R�[řv�x�	�l�x�����(�aR�ar�USo���_<I������=�$ru>��`خ~л��f��� d2$n���VS��_��y�\}�eJ4'?�	N|��h�ܔ�C��!:65k-/s�2�%�
�O��#�P��]��U.=�S�_�I�s��m��G�࣏0A1'�LQ"�b<�W�e��q���X+�E�%U~����ܟ�k����X��Y�y�GJ��]���X�B��P��)����i�>!Q!M��c�T�k�%!Җ0��\����rϟ�%�~%����_�u��!�'��%��_�Z!a�GY��Jf�*A������O8z�&�����y��663�pd2hP���^���o�`���A3�]�L��J��	��i�qWw��կ��y�=���&��{�K��^߼��o����ϴ&G���%��P�K�$Y�D"*gL)u�I_-ӓH+^S��ۇ�b����`J��b�?5��;8�{���ꢕ`�W�)JliV�V��~�1c�}�Q�t�����N-x����j�>乪u'g��r�6�9aC�0<��y1c6�q�3�~�G�	(p�����x���AD�o�w%�xq60V�$�l��A{�*["e8+V�q�t��fǎQ" Q-����J�"��o�X���=s;�0s�
�m�c8p�p�����=�[�L����N��;C�B���F�ޣSΠ�J��b�@H����0�����6��{��ɔ��}����/��o��p��*�]��S�P�-H��cO[�lt)�bo�>���R����q�H��5�jH)ɜ�k(�Y*�I����|���o2�-M��@���w:{'g{�$�l�7�~�7�z��Ì�tZ"��R�9	�f�]�#I2�`�����q���4r���W^�՟>���C�����Z��CH�*Yw�B��f/a�9�6H��82I�3��3r����s�Ir����4���~�x��U�?H���N�>0�I�L�������(m]U/8ٰ    IDAT�t�TJ8�+1����ʦ�aL�uҒ����_�E�\����^��������۪�
�� �y�=
Z�uP�XI h�'�E��[���g(MѨ�����J���:�q�4Ƨ�2�L�����uYI����jMp��S��^T&���T��U���:��{��v|f��9�A���J�` ��]����(f@��q�iY2�)·t����ş�%��;`�h\p��cM�5����j���
o����Vd��c&&X9gv�F�)j���]�p�c��sK�
�5�ڣ��B�*?Z�ΞX7�iRN��݅[�z<1�y	r�(L'�5�ȷ��`���;�>�}���ß�,7>�E2s%%��g�z&Y�7�s���$	"�3 ��$G��TJ��~J�1d"K����y���pw�2�d��G����O�W��qt#E��D�Ȇ�-Þ�6f]o�٨2%U)	l6�L�d;R��m5m��daC�6T��c�C�^�A}��z�Z^V-۞�:8����
!�Ԝ]�������]�s癥��HF3����)�Z�Cpgl`�;����8��	���C���%�QF9����`x�'�(6�}��}��?����1�)��B�����@{�G��Aa#�#�\ ��g3�$ޒ�-N}����:~w���W�1J��2�#�hi�J��{��'�ևk�f����{�t�i�y�R��Xl�xs�1)W؀7�6��@�%�`�Y�)O�s�2��R���	��ń)6���eGSu��Y����I�M��\� o�87>��0/1?��/=�V6@�%��ز@z�H��&*E�)�w��`�Q���L��N����q*Y�}k.�S�4L��iȋa,���V(��*hǢ��@D������F�8��0.̃�a-�`�rIp:�c)'� \Z�q��U��X�����	��R����-,��"�N�B�~����l]ά�lV_��A
����K����L����fdG�`GC���6���f���z�p�K:�_��XU���
!lR_y���})y>�7�O��5�`�Y0V��kZ���}��b|52�8s�x繧y󩟒S�=�ѳwp%M�:a0�h�p�"���I-qw��#�UZ��ǲ!W��o}習L�I�����_��$����Ɗ�r��t�ti������u�Z0��զ1A�"��{��>�J��{��u��q����4mq�G�(ޣ�T����8��-�N��ƕ��S��������'�A�{�s��9\��qx������mN*\@J��8���l0ff$��{������l�K����~�c��������h��e��u�[W���Q�n����i���"g>��W:��Mn{�]w�,���:G������I)1>�X�R��6��[ծUZ���w���[��[o䦏܆�<����� Aj���k}��>���j=c�{���O[Ч�Zׯ>MD�9n�-B�}H��D[�㽯$�~B_�� ^�Z��P��C�{lG�QK1`�$�z�G/�V�8�ߢ7_On��	ǆc�J����ԍ����$Ho��{u_���[��]sl��[��q�x�ެ�R	��wy��?�����t���1�Y6��^BQ?�[*wLj]�X���Mٝ���6:4Ğ{���"�]���{?�����1ز@Q ��'
#��8��c�W�%�	f�g�y_:�{��^��?1ȧL6qߟ�n�ܗ�@�)�b4N�N�d��+cq��\n]�[���^���ȯ�_��A�t�q��j���~6ϱ�4˸�w�gS��r�!n�������}��r�����w�	/��`ꘗ���y"�ԁ�W���&o&N�5�}�Q7����oغ�,�]`���S���TAz��NW�5K�o1�l�kq����;��ds4�$#�C�q����-�P�����S��{���
�-��V����1#������#R}��o��������Mؔ���r�S[[-b��g��0�a~���~?������{v��鶃���1���d�y#{'*�*��2�� �kc���b���:�Y$��T��keC0�K���v k	2�����ck�Ԍ����S��P�}J��[G�������x�؀\U�l	�G�,@h���p�׬[$���6¢;6R���(3%I�r;G�H���$ջeF�Z|�_Q5�%�1�Cd��Rx�H�}��o��c|�=|�k��Cw=��P�u$R8l]��R���e�$�F`-���#�E_}����>��O`��lpח���/�%W�!b"�i�0j���#�]�)�jlN,e>\	��>�g ��?�u}j�����_�u>1���)�(�(�gi2�j��:8�_�:7|�Ç{$���׾�-�lʑC���O(M;O��&N �E�z����t��)n���8��Z������4׋!���7+WL����.�ۅU}�b)��﹫��|O��L�+nH�y�$�L.��[��rR0�����Z��sjϺ\E���Z���;�Ռw���0�8�:r�m��-��٤q���>&�uX�B�
	v���k���^�}e�pt�V	�1��JP��-��W8��pR�ta���c��oIe-�P������~��R]'U�'�V�84!�����nWUں�ʍ�\�5Т`��7��T�\w�=�������®v-�쾿O��~��vLh{\A]��� G�w�y�U��}ңǸ��1ܼ3ɗC��r��M�2bK�v��G����T+&�͋���ŋ�H6���g����F9p�A:P6����H��5Ƅ�a:e�
v�>��`�2��翣|���bo��3_�+N=��\.S
��MZ��sDZR}F������Px�|ֹ���Ή���6�\�C��-n}�E|�D�Kл�t�:�B�f�[��)��̟~�[>�(�w��+d/������|�}홚3���e������6{qr��GN�y�=�M��\�՟���^|	��Y��/Z5_ eH�܂K��>&o��U����21>�>����3-'n��Ŝ��w)��$>H�އ"b�E*��+L1]ͪ��!�K�G����Z��,s5�̆�,��Ɛ,QX���E�v���Ѭ+�q_��ω��W���z����b���=��w�@����貃�!�\�Ң�$P���ZJ��n(~Y��cn���bi?#\�X}D��X8���7�o۠�{��E�X��W��a�}�x�I�|�%���J���#�G���&�"�����6��8������
�Xk���[���⶯"ӌ�����L
�l���{�r�y���X�j�����kg�-P�(p�����+?���I��-w0;~��)r�%4�HH|p��]-�Gp��g�T3S�Iiy�}��������B�[n殯�G?�G�^��,������͞Yh,������R���H���5]ַ�W1��w�Q}�.�5�����6AI�̸�o9��ԗ����U6�ٚ\��/~�/�����_=�H��р��
Ȓ���5 ܅�!E�	VhΛ����+����d�"�{������3Pr����,�=m�q��:f���������r�Q3�J%�N0<y��=�%N��1�a��WȪ�dƘ�O�Ξ�{\O��.��oѺ�W<g�ո�!F������l����%�{;Ӭ�^���ս���w�#�}Z�X{�'�����4�2��	{�Ĳ���M-������NZ������o�!I.��⦈a��[Oh�	�� ���[�_���s��Z��l��>�Q��s���3�/_@�%S%���8�^h]�*�R-�ٸ�^����Y�����z��66q�)�_AO'x!)U���:&�2�n�X.#����Z+�c���{�M��A���
�8S��q�?¿�*#�H����<�?|�܃�	J�����>R�v��s�H+� ��4S�>L9������<�o�����fds��4���ˉ�>�^�n���y��5׷��������s��u�Խ�+��{F�����c,�Qf���8�����O�}�8��{��)���߳�ڳ;<&ߝ#���,cccD�=ϣ�/Bb�Fq�$NkJ��J��8��=�<~�ɻ���?��[�)͜Y/|��A3H��������}������nF��O�/�k�m�8u'��&;o�ƅ_?Mzi�P2�䯉�sh��٨z�*&�ö�}�H"g�*[YZ�7~���y'̦����L/_ qv��+gvqV����"�111�kV��V�/ܷ��規�'n�:B��Ή���;��FV{�ǃ��/erj��.��SuP�د-�Z_��8�vU�}RG��$��&)[I��r1��%�CF'�3�ԂKk������,�>w�Fq�c���|<'�]�[��Y�~o�s��N���|���{����{�J���=]� ��<{;�95P$��q���`Ͽ���a�җ9q��p'�{L%��e0�-&�J)����x����8�AE�rnn���_���0���h6�{�i�P�!F]��򜭶sv��c�j����+�P/,�K]��n][~��8L��.�����4Ϲ�S���{������
?���wv�}�Nn�[NI}J�W�t�q%^�W����>�X�F)�����M� �{�˿{
u�2���v"�fM��"�T[�4����|�W��ӅU��g�2af,�q�^��ۂ+��e��9�%)�� ���&t���uq�Amյ��k=�h�^"�x�lc���y.��&���ʼwݴ�ЎM��ʒ]�[����E��ʺ1w�w�V�Ψ���q�M+h8�3-�U��>���a6�T��PEU�����8R*��Qj��ᆂ8���N�q���l(cD�^b]ms�G*�.T���5),�AB�rR�Xrث��
�`Z��3��>x	/����9���0��z.�RJF��5없�D#ʂB�����M]��n�B��b���s"D����A*��H�^ ,L�F�Sfۯ�����n��1��G>���Q�2��d��&'Qi�}I�w��F�+��[;��G��9^�5��a\�3p�q��`+��
�/��\>c�yy���&�/=Ki������ǥç�`r�(�-���2�e����D����y�Ph��d�k4H�Of��eTR`�#JNl(�>�s�����w^`@Ib<��DGըj��E0��Y��ε����I�k�kT��1X��F�L@���a��)��TG�*X��ߵ�7�PU]�["�F�4�h�{�}�xN�F�����vj<�`z\%����㵢�DHp�b�����?�(���v�E~�\���y�im��9���?((	h�`�]ԕ��J��!)�qH�;b�͐唽b���M��1����9v~�]�w.3��J�Ik=S�u�S����b
���gZ�"v�%^I�M
�fO:��4C"-!��'����{�;tG>����^${���)�[�ܔ�����%�ڒ�NXA�4Z�%;z�o`��imW��P�Q�
{�䈢@9�s�F$C,�,�h~��8������E��eFn�/�Z
�t����D��#������v��Z+"�p��M3F�<�vN���o�B4L�V^h�� $�:��x�ph��h��	��U�J���Dk2�h��/���^��b]Q�A�KrWTR�N؈:7%�:�d)����SJ^�-˹�h���ƙ����ն	!i��$	R٪���6'x��^���=���c�8�������wq�=�`��;8~�F��/1�L&s@�dBiBF,[�w��K��8�������CQ��(#x�7����������Ü��n.��c(�9���$M�̧����AmU��[W�X\�۟Xx@JAaC��l�w~�4��u/��I�u��}���u�+��x�,��6��b�����G����n�h-�`K+�stQ��S���5�;���af�����\Ĉ���a��i����&��l��;�ht��>�S���X���c%�kj	S��ߕ,��¸�\�ڶn�ո�{�sK�����%��y�����w����w9~�4�2<Kvp�h:޷���Jq9l��v�p��	���S���W?������O8��g�f�{x�L�v�y�_Ӻ8u��h�Tj�wX�B�L�!8f%\���<�/����������!���Zi�h���S�s^���E�A�Lg&��X繐��qE9��}���L�wp�ÍE���m`�EK�������+��ܷ8�<���W�U�t_�,�@4�����/n��ZWAo�
]�;Zk�F�|ٛ�dٓ[6dq�C�`�m���};��j�\���y�D�	��7?�SK�͸���[a��>%$���S��ԯ9��p���k&&Ś�	�u�4l0c���f}�|O��uj��?M����{RdH��<��E�_~��w�A=�_�2�}�8�#�Z3�Ph�p~���%�R�COR�.a�~Al��� �R'֢S*��9���3Or喛|�˸�[���_f��6~�]N�9�L���R˾�ʸ�c?i���,��3߽L��O�@z3�.��A���[�1�՝p�F�Rw*J���āvR�>b��@
���1����UL�⽫M=��z��U��!/y�����KO`��p�6FCv.�lFk�����b���x�N�!�e4�L�w�#��'���Yr�g��o��;�5�΢J���C�܇�I���T����{�T���J�Q�9R	�)�ؔ��o��o���l��;.���y�<w���p��@����~;�f�VT��H�qBb��_Z�1p�4�}�17_O�L��As R_P�Ev�f5� h@Z�w�[�E.��!5{�fĄ����ba������5o+�.���ϭ�6벪E����xs��(C�X]������񠻎V}��py] �80�:XԎ��A�!hQ�h�Ғ�g8o�	����qBiMȐe	�b�R���a���UZ��}Amۨ�$(%�O��r�5s�	�+?�g�������n&9s{֣�d2���P�m<���[7�����[z�Jp�U ��rƐq�m���?b^~��l������/�9�=�s�R�"�oI��s��gH�B�HLWB��@(��(!(�g�<�@�<#_0ʧ$�"��@8t=����~��s��cz�]����w�԰�O�Z�
j�8"&�
�cԻ�ֶ�!�{NH�I5l�S���w���Kl(G�%H'BJٺV�yN�
��25���0��q����#�F	r�>�z���O5���iS[�w�~d�VR�FXu���cR�P>����K9�k�b�������e�
�/��(ߧ,���R����z+�]K���-60��%BxJ,�#g���/p��i��o���ϐZȆc�]%��SQȭ�_�(�ǺXw�$�a�E�l�j�������:c���}�����1���\'@6v_���#��S_[/������ԌF�@V����1,��jA��lj���;0��nmq�c�e�ֳ�z�(Ci)M�%�u���@��ٸZ}�qU��!�2��!)��W�c���l&)�4��|���)�8d����()W>�۟n������>[(��p%�W_��?���8cٺ�.n��WQ7����q6j
�H��Im_�H��Y��ʑ=R �w�=o���)���t�p��f�B�L�B;Ű�2����ڰ�s��*� �p+�hR.�u�u(�b��=���C����g.�"JG��3&�^(1*R�S����Á����`�/F�����q�2i���o�l�� ���0��f��7���\}�fN���Z�Z��c��v-�l]�ޑ�`*L� �3J2R�Aa���c��؃x3a��3l��c!��Y���U�����Z�����UZu���C�v��çP�r�y��RL�x�b]��9cq�0�r�������7�H��Wݯ�:ƌ���u�w��jO�<ϙN�8S��P����zy��b��b��v�U\�h��	����;��k��� � �%b<`.��q�7�f��7Q�d|���\.�I-BU��]��}}�N�j�Ze{�u�&�")�S%W.7�3N�v�}._fph�M�}�#w��Eo�Ì�A^�+��׵u���
    IDATZ��3�~ݸ��$J`�3���d@n=��li��'ȥ���W$)g?�87}��L��d����$$
�R��1/�$�p�hf�!���ҧ8/$(���A/��e������&�dt��]ҟG�~oWSg���`w�x�o��u�7_�J����)%Z��1��Ue��Di�#�d>��x�Ep�޷��}�����޳�nbn��~�+��f��1�w��_���9�L0+g�$i(4�����9�6}L�*\t \�D���T�gHgH��}��g���M�i�`�}^�ѷ)/�'������K�B,�����5��Zփ1��΀ēJVP��l�'I�r���E�-���U���zm�kz�F�=�V>����t��Z���������wv����f鋛�)Jd5���A�Ѻ�n�׿��/���y ��[����ܹٚ���˦�������h[ 2Er�mL��Ғ*M��7�4���^���B �Z��+���g|x�`:��o�$���'y�g?f2�&�l�~��!�'s���~wzp��/�g��UM��pN	�Ba�^bH%���|����M~�<��QN�\���v�CX1_u��'x��#5�	H��L�-J��$>8aYJ<J�k���(�E�ب� x'���*3P��^3r��$W�9
��W��;+����1���26����bA�}�����"��`(fs|��԰՗�Y�p͸񻥔X�h.gǸ��ͩ�>M�N�^��?�#�ϿȰ,Е?�ђ�%��8saL���C��C$W�'U��$�b���9��`t����~��l�v����;�3K^8�+WJ�u��n,���9"�a-�/u'F�C7r˧fxD��.nB�����S 
[���S���u~���m����y��U4f��;�D�{ @���Q�=}cs�5N|r��šV�T������Ѿ��/?跾M_��9}�o���s��}�����dHa�/����>�_}���U�e��w���SX/P�������4j�`����1���J1/
6�c��kr�e��|�-��g|�3{�����bV UJY�+|"=H*9����xkH��bVX�N0v&ƇR������s��a��o���|}�D���B����]W���\��[��B�(���=���Xci2����ǹnX�e�v:0�2}�6~_{�j�ǻ�d�LC���9C]1� �}3�G���}�f'!�):/�.G����Pf��B���(��J��S�h���P�#ʭ��Q��V���/���'~���S�����m["�`�_�VI����0qV�`���O'f��S����S���m��}�=>x���;�d#�u��W�k��h���>}B�e�W�ջ/LG�����𽨱gr�����{x
��(��}$��}X�}t��?�仇vf��y.ƹ��q��隵����3^}�ŉ�Z�7��RY�	i�M�4�F�s�e	�
��B��H��Up�@z������x���D�ҍu�4�8/H�S��9�+�
�\�P��>�j�*�)�p����5Ll�3�����
��}i=��&���ak�jT9'Y���Z���u�wf���!o���\�ٓ��$g����^�T���sd�:��R���x����w�1'CyU�k�fBh��L����/�T`=�·�%zD�C	��K����!����O�������oE)�5���CvS�wӦ M]��>�Ԝ��4F��QJ4���ۆ��6�p����X/�B���a��(=�,8�0�����dȑ���oq��o�tɑCg��K���gPf��s������$ =�ȩ%�E*��6\m�d^���+����ɐV�l�eY�!4f�-M�z�"Q)�J^�GiAS	�!�D��"�B������V����h�3IQe�rM,��E��k���JZ�;�u�}w��B�I�������jU���u��CkP:��� 쒄��J� G�ǭ�|/B�� �){0*Q�%�l"�Qv�)z���^����|�����S��>�������m�qƱo������ř�<�!�68���ոT�	t�zu���hT���BP�SX�K��b��a� ��A�M���"��}ʝ��}���R�lZ�&B�N"�lj1�w,���2TީցS��$h� ��7�k�`W���g9r�,���O~��l2@�e��D�EҘzMS`\��6�<��CK�l�<0����k
o��ֶz�JJg+�q8�ک�M�apI�����oq.0�R��Z��Tp�ᩄ$UF&^#΅PJ�@Y��M���t?d_�N�_#�{�^_���(�\���;�e����!�_6��D�������3dI�;�zA��7T���,I�LI�4�yl>g�
f��^���i��#������dY���M�VRs�Q�%���&�O�����JR"0�9fyIQV%l�A�&\|��*�(���z��̝�"�t�C���V�CWJ�^à�$����h��4��j�a�JJ�����p���{�)�d����b�ɇxS8.y�J:!q����?DH�-dP�_#qu��7�`�] ��{}>N(���|�c��f�k��V\ם�>8�!�%�Up뻯�7���Vy{l�V�8�f˔Lf�c���t�S�ob{��'�r��	�>� �c)歗9��? {�<[����/wzvny�I��Қ9�4����Z@�e(��tb1Ó���O����W^}�|�D+�V[4>M���>��Am����Y<�t�l��H�I�$/�s�)|If-��mfWv�ΦJ`3��Vb*!�@�bD���>��O]Xt���U}�\�������I�}���{�d�U�M��
����Z�ݭ��S��/���`���o��T*h�J�PIHc�@��%]eu��/�����$�9�Y���I1e�	|:�н��n>K���L"i�Yn���\z�e H����Ͱ8YԆ����wg�#%��Tei)M��J[��|����~��1l�� [�|�+zLi�Y��m���{��TO����8�����E���m�iˮ�#)㝫\���p���c�}�4w���8���q9� 'EZ���=��X�S�%���z,��]�^�tk��`��a�Ols}:�c,#��9�?�~[un��F�,z�#.ۼ�1�C�q���bl�6��c}�RJ��1�����o��?�}�S$�7(������#�~�}��S����:"������+鋊�ׄ�� /���M�(��������8~�Q�~�+����ؿt�$Q���<9�-ێjm�]�Q,��b������q
�B}�L�ds���/ɋ}4�y)�<}��w�Ed�$�"/� fs�T���%iT�]���fn��k�V1,}��6F���%�֛�`�<��Q>���b��g�k7I5]���a�g�º�!�_/��&���u;B(�{Jkp�C�9�Ϟ�$IF�Ɨ������9���:�wJC>��ʜ�^y�٫ϡ�����g�gv6�,
�ʌѷ��	K�F���֡�l�����'�G��늵.|1�@��IS0�9��_c��O�5�c䈣�s��l�\z&�f�&�vh��}�11QlesZ���UQ�����yCY�Q�LqH�2�y�9^�������>��y�v�����������,�ȵ��{�Uw,�zM!Z5����c��w�-�����׵���UHg�s�U
Z5�x�CPU�50X�D�C1E�g3�Ő�b@y�&���W8��/0�:���&o|�8���1��C&�K��>�sC��qe9k�I�ȯj�Ĭ��z�������:K�2���r���[�r���װ��"c�#�*�����X"�MDS'��Z��؈a'CC��,`s�;����r�Λ�3?�>�D#P�M���G{�0{׾_��t��p"�5�xNW��N�`&����8���W1����b�De�sU_G(��,ttQhe"�NxpU>�nE����>w	іqd��GoE�y�LQ2��2X�k�k�B�XV�.sh!������<��\x�y^�'��E|"��Qv1�Ō����0JGP'&Ye^lXIKU[;� �&S��\Y���aD��v޵��jn�dI��GgI��	{�?���.�o��O<N9�� Ȓm�M�=��qܝ�*�{W}]��c��W�$I0��W1o�{�\��6(f%���Y��Y���ߢ�N\ϝ�W�{�s;E(z�U��"y�X}��^K�-8x��V\%�w5��'	�%dS��ܥÈ�뵻n��_uni� �]W�3�������� �G�伮)Q�A�m��!��١��ȟ��?�i�7��*�������.ٕ�l�v�B�m\W��V�7G6����b�"�؋Z+(�/�w\�;Fg��/|���G�y�\����FZSZ�)C��n�u}�}���C��Q���H�h�a�(�d_���N2<��2����S��:M)��8���ЛZ���E��[��ץ,]E��c�����ܯ�<�ʺ�RF�5�S_��	�㦻�lk˖|k�H,:B� D��5���ڄX:�z����q�aƙ���G}��G!�!��Qf�9Zhyhvm��o�fr���2���ْ�ܛ���l��H5��psC>����b8
!��/�����^﵄������Büpg2��|�5^{����d�1�~����^���m�T\E<ֵ���s�.�X%��@��Z�r�!�Z�dB�?g�fX�4�2��3���o�Żob��ԃs�W�Fv�}\	Ji��/ES���^�x�\�A��wh�_���G}�)%Dk-z����R�A\��s�����>\p�:sU_K�~)��/|�>³f=�3���.�������O~���o$9�����7�Av�<[Z1��$^�)��7��Y^+���ܳ�3;��y�0�x��X�0%�sE��������%s.=�o>�k�tJH����l��5�s�M��mPD��m�BN���5��|(Т��y��[��g�:sz�1����+��.b��Z�����t�Ԏ���zL���w����d�a��s��_֚���u	|��-z�a[3j/��T��.�#��,�\T��hԹ��6��V;vx$ߒ�?,��>,9��/�1��Di���ҵ�$u���]��DdH�)�cnL�(���o?��é3��G?K1�7��*R#���.�0��e;�� �f��'X�xs�9u�!�%<ޕH	V�� � 1���'����d�3<s��>�i��[̬i��kU]ۋ{�����DT������j��}	ǵ�$�@!�D�0��Ô�l�,w�A�t.�����%��.��y�����3�O}�wsC����c��T����R��*u��aQ{��Ҭtۇ��W�>�+����h33ײ���a}�pk�d4�D,��tr�5�b�%�.a;=�u�~�[��ǈcc�r�x旼��`�ʋ���[��2V�&�UD���e��F=�.�RT��fVEy�d�<}'�mwaR��d��ERg�o��R�T��t�������PED�Z}�gCD����e�jt��b���3���C������l��E8ϦL�sp�_V����c_�Z�b��2s�ժ4�1�෪8\mF��߷���d�+��t9�>'�%d�����x�u�9Vhg�����jC)��>o��I~���s�Bzr\ N	!f,�&jI�b!Q�G$�$�e�PJv/��_=��J������l�:PJ2-����a��%�8)eS�O��"Ͼ��ǡu�S&� )1�N9�4�[o������'<�>��M�3�L�8�X�XN��m]g���|SkSt���ocJ���nk|�1̋)�VJ�g$��,���D�26M����+��'ʷ�5d�{9��@~��F�R�ա4�����Vק�[��X%�߻�X�s���>��E2�?QY������U�zU�[���/�`���p4"IӦ<�i���{�D��O��|�Hn<��S�{�_x���O�_��c8�8��[��L��ڱ��ۙWq���Z���#4��y1�@q�C����|�R�x��'x�?&�M)˒�ܠ�4�v���%�s_���5m�7c�����'ｇ��c��p�W����ʣ�Y�8�ـ��t�.�ר�kH����ݳ����k��v�W�^��*��y��&�d$d�m�[""#d��YY��
�O�B3�Ҍlsb�;��R/�x��)���S̩m���1��9U�s��)�bXʠ��!Mbȃ�˅�H�L�0)ɼd�dH� �Gy��F����hHjlP��G�<��sr?'�	I�tء��b�8��@2+Kf[Lo8˕Yɖt81��AB4&�:v9�% ���UM��!`5B����ⷢ��3I��x�q�D塘O��T�0��M��O=���'?�5.om�C��49J�7G.�����Y>"@֠$��m��I��͚Je�Z��&�@��ȌDI�R9j�W')����(���!������$Q�����^rx�W����?�G�7IT�������r2�+�U�%�,�+�qW\Q�	X� �&X�/W��>$Ũ��M�u�1�]��CQ�eY1�$ɐ:�� ���E�^�n�q�`K�H`>�Ըx���E~AJ�: �
��&��� fpʲd��+�w�q��Cׂv�x����}�H�L�4��2G����gN1޻����x��'��p��|J>w�J����n���0/@�H���{�x
B�Y[T)D��W�����X���"�dN����l���p�L�����-O�����!�\@��i��H2D:��?���cB��|���%$D�N$���:��J�^vN�
-�_h~��.;"%�6v��;��jy���O��P暡Q8m����p�ܔ@��5���^�8�#�A� �8_k	-R:�2�����,�u���@D���W�u�����M'z':9R���Ysv�����#����sf���j49"EQ$�Eшl�ͦ�n��ϻ2� ��DdD�k͠N��ʌ@ �����l�)�ŗ������!����dr����>+��ೣ
�6����1�3�|� F���}UU5I�]�>G��ې�s��|0�@��3VR�X�J�4Y���T�=#N5���؁8.��lLq���[��~F-t�}��9_���P�N�g��ֶ1������L:���"l��}>�~ظ
{�2/?���p�=p������'�V���`�!�5#���L�`�M��$E�$���#�:�~MG
��i����^�7��6���-�cv��d'�p��W���q.�]B;˙�.-�9tn{�A���G���߱s�t]:p}���K�"��E$���lF�8���~�J���P��.^a�R��C��%1����	A���G�t� l/3U����K���vC�u����.�}�Iׅr���$���/}�vƖ|#��~��6���޵��e�6�����S2QsNnYn����C.<�峯0ί�6u����hݮOO���QM$�
��f��k}9C�r�(�*���'��
��y�Z�]��(�<�fy��?��/�EEG��9V$��a� ql�=*���s�� m*g�\XNq��G�g��a/\�Z��N�q�Ca�k둔�m�Y�|�K���+O�T����/#x���i�Q��Q*a�=z@����O�y_�.�x����ݙ5�N!�+IC�]$��L�9�q>eaچ6cD�&�-��[!��26��x�iRF2���VB��1G�v�Mc��-M���W�⩯�������sӻ���N��Os��I��-D� S�5�p������ƈ��$��%��;��g�R�������a8s'��ܗx��Y.��,��9{���N����^�`�f�H��9��'��<R�!�i�f_�I[��)эO8��$Q �`e�9 c����g��/���o�̥��9�Y�@rf;�j����Jl|�k�(x�UJ�Qj�f�
��_�t���y.I����D��1�C�0�H<6�!X�H���i����U��ZdLG�����NB}&    IDAT��T{�\|�)v�q�*^~�I�_����TY�3�&�N�]�mk}Cc��4�&v_�K��й�p5�R�R.�k��Юb&�}���}r�g����i���s��'x��83�b�D8�����D��ù2:����e��R1QVv(������{Lo����/�����r�$W�ge)���y#����h��2�M��4L6
�*m"��t ׺��#�n�]�8�����ZD:о��^��8���#�g��������s(���s^����4�CL4V%Z0�T�'%�c�w�(�����\�7�(�9��{������E�F��>ǔ��o~�>�2�>�֭���'������>U0>9��kB�4Ɩ�2���5����$�t4}���TC�D�,��Sؾv��?z��|�C�Ż?�y�|���*�
J������1����x��͊B��hp��P'^�Ү�(9#�~>��]�S��[Huȶ8&u���[�'̬F�
�GƎ�P
����Ѥ��C���F�k��An�������J�0Y߇�z�Rm2+Xנ^�]�`��kk��Q�v#���Ϗb�iI������������/��{��\�q�O��#~sx��l���0="�4�R�3�)a��`���c�*h�Ⓦ�ܒ�(X���I��s��GXV�T��y����>2�	�U�t���9�Xȏ�g�?k�;��̐ l�E�)���N0��n��)�g������k&Y���]Y��"�#T����H��g��@��4i�m�I�s�L_����^��+��� ��xKb����y�`](\L�
Jn�%����˅gT�]����R]�"jb�f��tr��u��u��Lb�q#�A��5��p�
0)B�M�c��J{��������by�k/����`Rp߇>���p��A�H9;郓��7[c����C4�'k1sD��P�I^pv�*���O�7��W��}�UE5�s�ou�VK�hT1�䞙ͬ"Ɨ��ٚ�]��.�Nצ?G���j�ϰD��_����c��)\P.J��l��!��U�yx�3�}idh�$��Q
'�.4�	V�8�x��9���O%��7"� ſ;�9��KF�a��PG�hc{=�c�z�5��c�9���Z?7A�߇#�t��U��3�T��*�l�cW:ek�Y��Sq��~ƾ~k�i[d1�E�`# ;%T΢T�Y˄cr�z�{�F�5{�<ϯ��U����X�U3��_�X���F�P��M����k�Z��f�>�v^�V��o���r����M�5^ ✯b[��@���!7}C�h�M�_K��Թ`E�����0N�m<�w�񇃮/�>�9��M��qJ��+(43�\�7�g*7bz�xb��G�fp�~ƬCJ�>n�!�>�7����z�p���̵K���Nu�U�
G5�e~�{����ZW��u�a�ED;�J*�gSKM���f�	�S�H!,2��
}�/~�/����S5�����9g'����� �E�;M�����Z�i���0�#i:���?>�SĵEr�nι��|]�l�5�Rۊ�i�|g�R4�a���rJ,LZ�M!d�o���U��I�4��!�ٔ�tJ��>߹�L�Υټ�c�RkB_�C��!����	[H��!-���x�f��sC}��Pd��K?K��T��_�_���ݱ��;���%�Ղ�z+�L��p��w�"�.#�D���w�Ʒ]�T��jx�� 2�h�Fؗ9���㮏�ݓǐ��,~�W~�4(C]Vށ�G�%k��Q?c����5�y���*�Y���x䳟a>��x�e���i2�l�GC���0D��p�#� h)�g�ch���4)����������k�U�,�e����+�F%��M5���#R�Hg�}|t�l(}b:��gC�dk��um7�}����x�m�9�T�����2*�a��~�w�y�V�ʇ�H�>2�d�x7��?�F8#��N�=����}�g�a{�3)2��pl:c�7O��O��®XZx�����}�+��3r���L��Y޺�F��4vV�Ck�_��}���Q
Mh����T%��UeJ�6艣��
���2���D|RJA�#3�|L�éL7�<�i�<�s}'ʸ���ٟ{&����Z���m/	Ԙ�ۇ��w��.n������Q�L�1«\ŢZ���t����VˊY1i�|g��FF��#��!�#U&�`:(��SYJa�4ӔFq�{'?�y��ԇ��r_|���|���P�2�eL�d-!Ә��t�q���0�G�7t��=Ԝ@�������wr�޻��{\z�g\|�׸PT*
(}e��a������ś,��@�\��;�8�[Y����ӧz�Bu���c	H��BP W\U{f?�n{�6h�)�� ��Hs�	>�6J�nl���7����ߗ~[	���챓O٩/��\}�y��.g{/����kxX�O�0��1���q�nҞ�7>3)f,�\�.KL���)jξ��/��l2��c������ֻ8�;��|�։]�ǟ�Ci<hg�:J�m��ycB�Τ5�ε���]�5��}�f�5�ٱm$�"7��\@W�l�}fk리��&MG��[k}iek?
MH���F����Z�qm={� hb��t�*I�a��m}��3����~_cL}H8O[*8�4)�1>3�e-sC~l�R����WQ��iǁ]u4��x�sxGf����}Z/�u��g��Ǎ����y%{�4�~�S�S��o��#��4�Zpi�`6�byp8�ه� }t�
��#�e����9ř��v�䦆��p�HA3��ѧ���t E�󰴸4,|�:�v��>]+6Y��u��q�}?�?Uy$���H�,OH�k�B�5ԕO�b�-���Is&	K$fue1�`�7)�/�)D�d8�Qֆ�
D�Z2ڂr.�(>9����uM��^�*Ė׶M�����g|�4��l����\�1<ڍ�H�М�D�Z�5��K�	Ǖbo��r���6r�<������?���QhCb3ȝ�ښRJf�	����Y_v2�q芺�þ�0~ݔd�Z(W����Ø���M�J*��kC1�!+K
���;��������z�e.[ǩ�|�;?�i���ej�m]aı�k,��VT��Ρ\�b��%'��_3Y���V��:��?�A<��:�	�	b���,�(2��>v=��2��� ��eB�2�U�d2�21v��R��u�,P�f�gL3��W���o�\��%�\�pN0��D���Oʃ���V%�,���CkE�g�����\(H�N�:��	Ɵ��J���j�@f���#9�0�8�ߘ
h�1��<��Be���:�(j���L \��(��*�B�&8
�"O�0�g������#t�F-j�Z�Ӝ�܂��L`�Ju|V��T[!n�ut�J�ۘ69j��N��B.j��SB-�@�_���;���KNk�_S�2�d:�q��Rm���8s۽��+������w�*ٚO����"s�(��q���)�m�X':#W��p�A�������uM^��gS�G�#�-,
_�aw!�+��Qg��>ȃ��2��
��q�Or<�P�cd��c� X� �`��8�gТl�`(rx8�������&�������n��i�.�4֟M���L���e"P�'X�  y���$���r�)2M�b�g�d����X�Ϝ�N��SNp�VC�ˌ�h�N�B?�B�:R�{��$~?作�3��o�r�6���5���7$ُ��Z�bq�S�,wLUͥ��^9�l���ч9���9@y�C�'�L(�1v�͝M�g��Wja���8cB���9
k
�`���s��1�9fy�K��9����].)]�ɇ&��n����ס�4Z���)2jg�n�$����P,�4��4�^�n��Y��6$�&�ڂq3W_�(5�EI���D|v��Mp�o�m�1��kɰ�DJ��4A�E�+~���\�<�.��0���?��k�Z�y�5�s=3��4��G����ZS.�	fy�V��:��sG���;���;���g壧)��H�|l6�hc�-8����G�<�l�=A�
{P#v���$٣���%�����2g��5���BgT��Šzc[�N�� 7vu�ك)��U��M��D#�̬!��Z)V3G=�V7?�;7��];��|���IU�,ۈ�!xe�=���*1��o��c��߷Υ�9u���"�h���F�`��4Β�&�y���0z��n8Y� C�J%�5�-@���nhrC�9�}�gl�����̱?���
F�Z�I��Q5���'�ŕ_�W"�NR��0�+O��&FS{���9���aYG)�x�l�m�T;>'�-�gc�NS׊�$C����g������V�1y��������b��(�v�<�
ɍjV2*k��
Ԫ��C�Oa��>�O?sVc��{���`WB�����5;�>��hj�����֮Ɋ��7���3߭%iR���ݨ��2�QU^�H����9ua$͕�'L6�!-h����v���g�s�kJ,+�������sC�8�%~}�0�?#���K7�M�4~#s{W�_�)�<ck�$�9�}�����L��ru�k�|�˿~�Z��V�Of!�|=��J�wð��mHp�7��2 6½([3škE���U!�ܜ������CԹc^���E��"'ӹ�O=X���Rj�b�)>ƴ���,^�z�Xw�Z�>\��b��x"��Q�X���:]�B�A���bl�UB6��ϧ>\�Z�1}��h�h=����
��#	� �"8i��V���u��amC̽��3�A���R���*�t�s�W_���_���C�s��?���"Y��JM]VLD�'ݰ����M��\Y�0]w�ki��k43�ZAU.��
WvY2����	��k���oQ����?���{�����rЙC��K�V��'��=��i����~<�ǰ�����m2W���F�C(l��1ږizA��q�--�\����E��͙�+e��Ic�wƟW:��	>�|Sx�}�=7ʸ6	@Cc턲,)˒LkʲD�9�n=��[Π'�Z��M�~6�(DX���c�����/�#�
f��g��݉O%�I�]�_���)�b�Y�u�5��{?ĭ�}UR?�S^���Bv�,;��W5�P��f�n�q�͵�yߟҚ�Գ܉h��}(�͘Mf+�8�m��?����f�����_��^`;S�Y�\7�ni��8޾7����m0��6eZ�5�oe��7L<�?>�	���'�uR���jL8b�G��=��hQ>48�ɋ	d9Fh��T7DE55{ہv�/��π�Q-ո����$7}��/l�	!�J�L{E��|!QA]y��Za>��θ��OY��"R������Zsx�d6͘N-T�r`�#�,;ڞZ��M��6�/�c1�jq������\}��\������'�������~�7�U,��e��P(��B��dz�PWל���M?dn�v׳�o���p��~}��٘�)��֕��j����q�}Bt#�JC�dL�XBe�������w�ocK���)__��,�˪��
��c�٘P.��w�7�@�pn���IK�e0#�D�0�����n�����f��59g�0}��{��0�z�7������/ٱ��@�QU����������x���k���O��.�3��l�}Xo�^f
��W]Bm'���n��b�����7�����^�*��ۻ�(w)L������ ��?��=��m�KkK�Y�S�����Z�{/���p��!��]�0�L(�"��_3��w:d�Z7ʹD�=;B�!��X1���h�Z�f��hUUyM���I���c5�|F�rTF��9^�����4�Ţd��G��z7�L��Y��Bl�E|��P�_
+�3�V��_ւ�wޟc<�o�X��R��{��q�02g��
G�{��2��vNy�,/��WY��g�Ɲ9���'���:���47�2��^
u�|$�h��Qw��ک��3�F�u�X�%e��ŵ�m�����Q7�F�9�
V1C�R��]�Tk̼Yi��R�0FXS&���1-w���t�Mߥ�;�wk�M�(�����k��m̪l�����104�����?gn}�����3��DF�]I�/�坛uHi<�����Pc�6��� �}��������.��\����E��:�s��IQt|<�8����a�\6��5�޵γk��;�`ɨ%êQP��jr��Gc��[�V�Po<��86�3ۚ3�LؚL�"��0.<��1&8'K'�sB]����1+r���o��c�fc{���Y��ڨ�Ǿ�a���J�+AQ��fY6��Y�Ov�c��d��8�w�e})$��K#�:���E�l&ۤ��x�ŏ�N�k�"�4ٖX���K}C����A+���vd�b�\z���ٳLn��[�c\�.�����,VU8&�g'X�|�<�M\t�a$����8��9�l#�sh��Y�5X�P��3jq�L3�r���ᵯ	��tN�ɝ�m��ǋ_��Y]{c+)P��v���P!k딎aӺ=���΍���ڑA�6bֶ묔jM��=���5��
���W�s��	����\ȃm��Xˡ�}��^��a�:�1I�yzdӌdTc�cZo�_���Պ|Rxa�824�d�萢7���Wk�����6/.�ũfC�����$�a��f=Lاi�Ԉ/��0�1�Ƙ������ʾ#{����9�[`2�⳼��`��ŌzKR�"�H��
�v��y��[e��q-�%�;�;gP��w��&�%�(t�S�aQ8��ʛ����|�3w��|Ỽ��Y^8Ǵ����F��s���;e},��ioZ!�;:�Mi����n��l��G����c�/OW:�B�.�`=h0عf������ lR��r9[C�P֧U�8T_{����	�R�	3��K���yHR�!9�w��__�ۄ�k�;�~>�B�rq>�b����Z���ckK�������mV�K��	�w�79��SfǷ�,����6�������3���hSӦ1�ƘƂᵆ��5��TՊ�5TNػx��V�������_=���j�8w����ATqc}h�$���힖a�wܜ����+2�x��ZV)�҂����""d�&+4�$c2ɛ��>%�����6��,��gc��P+�M�-Q��P�\�?�&�3�?wS����}����~�$�i#�DHi��f~Ƒ;�$���z�c�{LS�ǡ���Cs����h���G�CsK��k�i-"��ﺗ[>�i�=�~�3gx�����_��_?��_��H������=�
SW�c�k�c�{ֲ�%嗵H���JJ��(�F�e9�\��T�Oq��q�8d��׹��s�!�V&hr\E��ɟ/Ҥ�f��5M}�Rg����W�ﲮ(˲ɑ1�q�����u2��$^�]���W�з�q�>M��Ve	�͌@�߼��k�����Lk�$?+�\��ڪ	qd9d9���%�D�TcW����ΑiE�Z	��@m�����P����Ө̠s����p-���(P�5Ue@it����m����,�3�n��C���Hm�V�Q)��2X�i��E�c'�(f��/q�s�PSn��>.^��OqKU2UV3Q+�����ْ,"���%��@D3�
�����Y5�q�L�Мr�ذc�R���2�;�(�G��V�4dK���������;Ǩ�.�ۗy��W�:DdI^.;�Ńǵ`�Iȋ�M,�*(�՜�P�kӸ*�e8�kc�E���Ƅ08ʅ��c@J+���U���Gy��a�k!2���葬�Bi�xk��/�p���њ��<�B�Fg�,�}�h��@��4b�c�vX#��m��/�,Lm�ʖHE"1$�FFM�̭s����� kE�k1��.*��8A�y�	����y�9�F�!j@~�[��X�X����$�J��HS>D�����ׄ�xf������i��s����ёH�Ǖh	����E,[҂    IDATY�\��Z��<��U�J��	b�q���]���C|���5��-����^����	���35�վ�8�D�G��ΛL/´ŉ�!9ŧTh����{���Zh��UԜ����s�YQ_-�Ώ���_s��L_��_ǽ�<RW��Ǟc���#�h���R�:��5�վ��rM`o�w�#�X�qHg��.�:�T�,/0�Rc1�0�t���pz�`b���V�0E.�J9��ʆ<�VG�+�/gq|x���4��(�YEchvItU� �-�1�#���ߏ5U{F?$�������(e�D��OƵ�w�����kH���̦�Zq �.�vt#Mōe�6�u������=����L����ݏ����;���X�+��2jV	N+$��o��pB�_~Mx��US�� }�b �֙����-\;8$�Oɔ���sO����E���я|���_�:q�l���\pz��!j}l1n���K�u�[�=�HHǖ�����9E��O<�3&y<]=ShC���^h��6� ;�/l7렸4���e>��r��7u���c^��a�%l�v����~^���Mr���W���1ؐU.��Ɲ>�%�9k�#�}z�ZC��5x��n�.��3f���kB�H�)���-p��,r1��R�`v�ny�}TԜ�Ѭ�x�7~�E>�0�+�ѧ%����ҿ�1�m-c�m�S6��2�&,qJc�NPm�ĉ{��{�!�*^���W?�!���L�W2�)����c��t��x�O�c�����4�v��wS�ԫ�o5�a´�e�����<�黺<�K/�,V���v�-�Rqs��&͖5���[0_L`�0lF�7�f\��(Di%��(b�r	3i?;��H��ݮ�B;P��V%��>o���p��g��ӻ�����p� '@ؿ��ju#�Љ��&|fBߥQ�	�_ǡ��{UcR�'
QJuj��C�t^���R9��K.~�;��w_��/P��}��'���¥|�+�0�![VLvOx��xӷ�N��R�5�1��퀺���y��H�C���������t�D@pު�׎��sA[i�E�ͨ�:�h�y]��zm/��x�m�C�uN�~�������yloѡ���t�B���fl�O����0�\���%��+؍�(mk�z���9Vg� �d\.�\���]����ԧ�OiʃWy�{���ϟ帚0��ctㄿ|�2F��m���xR��s.��V!����A����竜�-�q�����%��/b._b�s����*�fX�c~��n�s�M���k�!�fYA�,�r�ZTL�B�Ey�:_ds�ɱ񷏷�]�;���^l�a�p�	Y���N:*�G�X`>c�ט4�^~�ZF0���z����5��8�Ƨ��C���싿�7��&��.P�:ͣ_�#�[倫�\�PV5��������Cĳ��+�E�|0�)՜�E�("m�������|F�*�
n>�Cv����7x󉿥�r�;���c��ܗ9?;Ƶ�a���g��J�����Wc���}(<���7��Я��C��p9׉E���[�����!�Y����m�F��Z�kۄ��!���D�Ƙ�&��F��fa~�]Cc��0��/��{��Sgl=|M��f�w�����hi��
�W��:eNCZX�5[�ǩW5��YU���4�>����/�|�2���_��w�`V�L�������$rQ��D�˛���=}\I��ZMhjl�&3d�D��+�z�����(�˿x��g�e�,�u,J��'�25��Xǘ �*��o��G}����f:�l�S�z�Be�l:!96�4Cvw��<�Q�La�~�����]�S��IDQ�pN�����F����z�G��� �$���O^��3�{ߍ4A9	grґ�U�����I��g�����F�sΟ��N�t�?G7ׯ�����E8u'�{�{>�Y޾zs��L�XGFP�c�@o}L=3�9�uӼH�j��a��g ��dV�����Ĉa6�µ���_�����S�O����1���_��� �	�0^���U����g&�\$&�ǭ���z���9����`0�ڧ�m�����[�1�oC���?3v�5�@�I�$!�k���uPk��%��=�n�jcL��}���������;�=����l��i]H����E|�q�Bu���^CZ��O��qhDM���e�H�����86�Cp����:^������e�����L���t��n��?�I���_���q�α��,��u���ww80���s׵Y�a�֎k�C��W�6	�@S�U����l��Q����z��������]��w�͕�<Ǥ�52��󌕫�X���I�ӹ��o#�R*$��"�����C��^h�3�	�5��o��Ϝ��s���p���]�27tgh�>�!�B��K!�4�w
���hёHmB0$y��I[GB�}�/�86���y�@��3͉�}w`�1����F3�y2/a��:ɿ�N�gu�M^x�p�L&�y�)��Ɓ̉���"��\p��ո��bmV<�M�M�P�|\� �cO&�)0�ú�T�ܔ��]�ٯ�{�=ԵK�7�����S��B�Ga�XQ��x֡���qN�ZK!�\8wWm��RɺV�"����e��/�qԵ���>g15m4���^M���3��>�Q��(�c��6�M�k�����bӻ"��#e�}24��wO{��}*��[W(�l��<����\��c�ZYU���b:?ε���{��c�ޛ�v��WƫO|����8��8Xy���:�O���oԛ�m��o!��]k���v5z��u��������>N��ٗ(�|�i�|��"G�
l�1ٴ���J�?�ӯ��dl� ����so~�.�⑌�c:��9EU��
�L�	f���������^�HP��.�<��i���`���
p��8A2�f�t�G�#�$JY�;�Z�! `Z&����$�.P���ͳ2�����Y*�s�lMi�Xe9����3O�ؿ���r�G?�խ���Wߋg����Ų�#�7��+&����""D��Y� $^p��%�4�@��Pe��&F���,����cs�/�΋��do�J�*��w~��l���?Xa��U����ihӵ:�[K%BM?���Ou�}|.�!��PjW�8�Ņ;����/\��Wt�c{J�f����1�z�1͔Цi����}��%�w����h�.e��(A?M�}S�Ji�����`4�	Y����^B���<�o��G�-�,Ϙlg\�+.�SL�-�{o�./��������q�����%s5S`�ͻ���1��6y��Z��b������9�nzN��˹F��ӷR�~�o>Mv�M���_s��癉f�ZQ�5�\��*��<�
"c|g/�|T:4��O��x���������(��)d��{��{�ư�(Vdx�M��Z/����6���x%3І!�l��y��R�$x#˘T�~�I�N�SF1<�u`7}7�s�h�#8(�8�).W�-��/^�K�ȵb9)��#���t#
�3�"`���5	8bB��>��u�O�Rc?@��$�U�d�j\��X��W`�k���1��ϟ��'��w���]n~�Q���:s;���G�*�P�� ��m�Tc�`��k]��#�t�ڽ��_�#V� 5�*sd�����_�,
SCڴm<�d�����i9�~�g{���~�H�D���ƈ����[�@ژ����1X m��;�����Z�Vdݚ0�|�W�4��+Պ3�� ���غ�&��%�|�\�ַ�r+��q��)�	�v\������r�
Y�9ƪ��u()����_�?�(`ge�u�y���͏�����z����E�3��Bx��BI��bI��yƘ�&�O���2�5ĜS�1����|Y��`1��
�w��A��Y�&�Ǘ�+��l�Z,�QfQa7�����ۣ��[}�O�ςF��&Dy'$�|A__��ly��d�PV��Z�'��$-S{�j�6Y����߅I�3�
T�׎QSm�T��18�D�D���2�q>vT�����3��Ћ��S�>��g]��ו����W�'k-Z���$dL�WrB��*�N�ˊ˗^FMrn��Q���{O���a��s�.���fS�5�[s]A�@C����nu]��C� 5`�n�O۰E��Aa�:?� �t���������jJ�ԙ�ǹ\g&s��>�.���Rغ��:y�c7����y��Kc�l�p�c�K\]1Q�!��v?����0�&�:�;\���m`��F������pA,Jm[	�_
<�&:F=�y�3�M��҇;��\��С~|�k�7\8Q��:&&J���ͺ�3�nb��r=�_�W�ȲI�.�s���k���9�$KjL�)��N;4�5R�%��i�?�;b�l�
�������ՇIW��{5��h�)1�'Il���}0`n�(�|�K�Θ��p�ykb��4�`�C	T-(����V��v�\����/q���?tY�׿����������h�"�R)��B��ϳ�b��k�e�RhGK�1���cB�� �5a�,����Rv9Ԋ]{���c�/�O����~�kO~��3O#u�Q�4�
9T��lN��T!,V��`@`N�Y��Q��b�X�K��ujQ���A	d�m�W��ղ�.N�v����92#L$�hŁ�,�3Ϫ �YG.��v ���Z�`��[e!�X�vhmP|�b1.�	ˢƸ�+{�n����F�P�澔�E��}����ퟅ�p��0Ԇ��J�����{��t�Q�����	"����m~��
�l����y���y��%�����ũ�beg�I�U������eI�,;��5��x�A�M\�N�co�u�SN�t��k�O������?�z�nYVh�x�������$C�5��h5'��r���ޙ�c�^(X$.�q��&�1�X�����$Wi»��~Y�kp��φ���6ͦ��𖀡ȃn�~���W��'6�l�Zm�$;�q����t�c�=�|.�5�T�흴!<�7�;C�}O���%�K�����v�
d�@�ɒy>�P[��7C�{����/s���å�\��S����w��Z�x���g�2��j�y߻�1q�r04�� )�����,���l�6�q�3�듟`z�	
Vԯ�����>����Ǚ����m)̚,�t�^�o(�J�6�����;��iq���w����j*-j2tc�<1@$;�I��I��k�ĈbC�bL�������	���S��g���Y�Q��ZY��7p�&�8yI�$���
�3f+���_sṧ�,��.�9v�#,�)R�l��-5L���c�cDoh^C}nzG|ư �5�Tƕ~�s��~�C��P<�(������a^Z.�����_��,�<J`d�ݐ����N}��O�˄�}���z6}OJL��t���=ݵ�5(�ڽ���������	�C�2�}��X�����̾=��&qR���[li��)���#���D�����C�l�|��r�`�����ȿ��)��%�k/��_�5��3�M�Mƌ��u+;�棁8�a����[lk�ʑ�d,TI��1s��}�{��s�a��c,Ͽ���?E]<Ǳ�)����q��<������N�o�p3�%��	.��Ǆҡ��1�y���eY�u�n��1[���W4(o�s�16�5���@tX�| l`���Bt���
ª����:}�ݔ���0�t<��crG0�8;�~A��}�y;��"�
�,�vvٻx�W��Ln�n{'����)������l��� �m=��J:2�!ؤk�_�a���3�Zi_+�֟`�d�٧�D�wg������{~����4�g��4��y�$3�AM|x4ޣ8�.��>0����1��ǘ%g���b�Y�J�f���g�B�OA7��0����,���3*��C<�`㜷Z��}���敶Q¬"L����N�(p�%2��~��g	�fP��`Q.�jE>-�+W�I��?�sN��^Vn�������8x�i��9F�ո��os���I��;�� ��C�@��nHp���7aYZ�iƎU���Os�]�G�v��Z�ڏ������+)�����w�c�}L��5=���HB�mhz���U6�֗�h�Khe�L��J)��kC�-u��Ąt�x���0L��eYF�~�ZG���:���z�>��!	��[;;����?�'Kr>Gg�y���K�Zk�D@ag��J�0;!�69�]�a�`�.�S��-)��I��	�e��Ρ\p��p�Ǹ�{�>Ql����wp����R���-��!�e�rt���w#G�k=M4S:�o#��A(S�����L�s�+��_��E>��۬�y}�����y�o��+O�-��ʊI>�2��߹��֧�켏u�"F�6<q��+�O�6��1省/05�㏿������)u�"՟[� �1@�y��wG��?ӣZ�1�
G�ŏљfl���o]ctL����g���HF�qt�U�\(����4F4�����x��{�=~yQ��/��W�?�|���� b9\��'}�4"E��a�2�����_�+�:�����*�Bt��-��(����s���v~�}���Y�=��ׯ0�&J���i5c�GDlRR�\�����ZS��H]�W�K�& !S� �$XK��
Siuݵ=�߂�Ĩ�KSO�H?Oߕ���p����΢z�����1�Ēz6[kq��FS�%2߆�'A:�!$�ZL_{�ݟ~M7�?wE�_T��;�N��'�}����'�����\�q\]	��	���s?�>w��Sn~�a���/rn����W8�������mW¦�Vc���gL88R8��m!ͫE^
��������_��/g��p��������������um��j����H�)���H']�27��w�b��Io��$-�S�i�m�������Je��ű4��k�ԯ��|��CM�}�-}��Xߩf��od��%��>�_�����~&�>QNi�;=JH��S�G��}z�Z�����eQ+��S���q��~��?�!��Ex�^��_p���ㄲ�ιv�@������c�#l�F�m�ѽ5ڢ��J�䅠ܔ���ř�y�3�ǩ�<Ė�̅����_��-)P�)ui`e���Ctip}GBK��l*�{;�!�xA&��6�2<b"�u�9� u�v.8��F���K��tc�\���Dm�� 4Lv}���Ûͽg>����e�㦤T����$*y&S���D|e��ǃ�P�	��3�W�k��dLjm��-�I���⿰,�fU���!c����"o����'���O���*�}��35+�&��1<�!���:̇^�90xf�_��9�a��V���7�a�p��O�-��<����Z��N���"'f\���Q^���|�9%��\L�Q��d3�M�<Uk�k�v��Νw:�L�g�O�G�쇄�!������g���`1r�Ws�ꆩG���c׈��$e\��هC�_�W)�<�����������_{k]����g|G���S�!著I���Y9��KX�v/����S��y�U�����w��s8�V��[ԇ��GҎ6����m��-�7:��?H{K)w�Ö�<ӬXrl�ѵpNg�=���<���W�ý�f�%�	a�Mp2A����؎y�r�����j�1*%j����a����؄����1,jǐ�7�	�m9��ۡaD�r����@�O̻�x�y�۵>�  tM�cE���}?����%�����#��xI�H�]�ˍ�V�[0����.�Թ���E͊
m���7����\�~��v�����n>����lM��e=�k�w�]:�>1�7�@�?O�*Jtf)�_�X6A3aoU2��تW��ķ�ɿ�?Y��,�-��{���Gq�t� :��V+�����44�M�",MU���U�����X$)V���U0�x4�����lِu����{u��0#��N`�%�C[?���!�;�ߐ@t
���j���_	    IDATyn�tܣ�����B`)�eٔ���^�L︝G�x��?���\<����7x���]���ڐO&���t'�1�\z�s��La-T}Z�~�y!A�M�Q�Pڐ�c�>� �mۨ�>O}����g(�"Wt�)˚W�FR��	��h�����oY�$;���(\t��*]�!<�W�~��8�Z��qd�r��5:/��ХҒ��$�L�1aA]� �ڊ�6�,cʼѼm�l�/����Oi�d���f�c�v^�RJ!�g��9��#G,���ڴ!g���FccpV��Q`�ҟlj���bQ!	�1����*ԖV8qDW�Xg�tA�"����i�>��� [g��5��uY%"�
�Ұz�^����������{�3��S��'�/������Ѯ��
$'�B��\���B�ه��GLB���ƿ'�S��c�L�¬�̂lR�����黼~�*�<��g>���8y�.g�-4�y��1�Z�$�T&����PN�~h��e~]�ʇ�eY���t��߫�sː�T�&��
�VA��L�&��y�j��5q�	��(���z_ ���ڄ � $艄�;D[DY�E�=��-A隧c�N�KǛ�ј��oDa�m�lk!�@�K�-�>׭���1��3�$濖u��pA��U�[?�W��G��@��G��X����I�rJ}�;?�g���?��\���O�������or�\�KVY�9p���xt��>��4��[k�ja��5��!f�ME����!Á����6��rb.dp�nN|ⷹ�ч��^���=�;��N�,ױY�������)�����u���!�V?�5�����lr�2�}�+���kqRD��k�܋�y��#F]8	V���
$�1�$��I��C�ZOw�����>�"�8�k:�?"E�D�����-�U��[�U��>ý�g��5�ZB�@f�Ap��;����
"����_����HB ��BRwK���v�ΰ�����9TV���+���=T�+הk0!�@�Y�8_�1�c����P�E��4����}f	 �{���
;bR4���fD)њ~�[�C��Xs�2��B I��$�%�P�kƪ��d�mbX\%+�Q�
�[�J��gU���>0�ZN��4����5o{}s�G�)n�ܾ��,軖æA���=�r`�x����v��$��wS�t�;�l�=��0H4�,�
��K���;޽~���	����"/@h#H���ӎ����E~�c��8�;�FL`R���g�Фi'+���`������_�ۓ����s}��/�o8Oc�<^T�(jb���I_��>?�}�L�������/.%B�l��ь�/��TS��|5�l	�Hgsq��e�̑W����(�o��9�����+���O|��?�Y��}�����J'SC�{.��.�;|7��r.�C4vV�����s&����� O����_�<~����/��7K��-E�6̫C{eQ��Ka�.Զ{4����
2=��08��50SF�Z+W�-�f��_Q{�����}u�1���=N�t80��b\V�)!�(��Za��X��T��A��BOBv7H�+oh��EN�!`�0�f�<?o�\�������8Us�6w�����ĉ������5����5���˷����x�/|�x�%NN^�Y*�JH�j��)�R����TҟJm���s��\QU��C�ʵeO��/����n�1����>�����Q�(��cI�)�/"�uP�y��.�c��;��D>�g7Rm��)-��3e���o̓�:F��yL�.xU�x�|6R�0sZ���}k4��>��^e��-� �s���:&�ވ��nƻ�+��Z�{��YMc�C�?�F������~☛��./��'�^�9��n�M�&��ߨkX������YNߕ��>����1T[a�pۜ�ڣ��=1��x�>H��#l�>˭O��>�w4�g���6����D�"0��Q쓋J��4��NҦ�0��ikPd�aե���D��2���(�)W�b����id�,���m� ,9�3��.�RF��Qj���5�&HTY��\����I��� 9���9J��01<�j�����	a�S֎�|�ƈ{l���6%�Y�L����B��RY?����?�]G��=�v��_����<���/��7�8A������c�}�t?��IES�~�����(b$.�}�
�Ê�U���-j,rP���6G�*�������RK�8����M��}��2Ե��5Ɯ��Ρ\��y��/��b
L��dO�]jטj��$m%	��<��>�B��[��Tz�eh�Ϧ�]��H�ͽ�V��$���1}_�̍��6u���������U�|*^�uT@��mMߟS�[^���y��b1�9ˣ%�Q�5x�$ؙ�u�p_��%�$0�v�~!�%f$�G1�ytq�����w����E��������>Fu�6K�TZߡ�BLP����!ND,���2�6��ӳm�$(�^+�ӕ%xj��XSJ~�1����&m��b���~i>�9a�����Ԙ�
. ��5N
�U|..�d���X\��Φv���D�G��D>��O9�YU�J��3|_J�Z�+�B���|6�`�YIr���a4�))�0��!�d�r�;^����ђW?�ל>��OѾ�M��C�ŧ�Fw��U� Zm����Z�&~��HO�73_�P��;�r�齉��t�7�=�����7�Su�]��h������Gb��{��!�@�S��4���3E�ss�[�dݞJ)Mϕi�۲��~�� ]����|��>������u�<S)�
��E�_��ynF����GR|���R��D��Po>��H��Z��+2DZ�H[������ �n���X4+:�,0��^�d��wI��V��x���k�1 �z
 ���!7Ϡ}�-��7�����^|�+l�}�kG���=j,^ޥ:W�t�"�>.��1#�~��w�aA����Չ�ԩ�ʥ�$��%9��+��)Ǣ�E�ke��Ąs0\e��b�Mo!�6��on���K!I�	�����o���Ez�@ħ�����~���9H^�w�!��e1�䧮c�;1 &�v�~�V��;w�s�CD�]��
�V�v ��p���/���?�#��ȣ4��Gt�#�� �~�K�g������o1�����#����͕}���Mi̗����.�ﰨitI�g�;G�[V����j������w�I�r�%��{��5���1�ٝg(&s�a,a]_\_��6dzJ�c��ȃ�ar�+��u��hj�]�Q�j2��͕�v�2���M%�9��v��z2�����Ź�f#vD�GUh�0��$d'���̠�>����z��RU�η��W1�(:1B��kC�r���\;�ʂ~]�v"H�k�d.-���k�-���'w��_�����9\:�]H�䍆h�N��c��bg�������jM�Z��v��n̨�ϩ�HW��o���m2WgQ���ݿ��D?'�%���s�^0��ڠf'Sc�?�#L��0W���������Ġr����d�nssHj,�\Q"��N��m�'H�y�lSv���8�J�xw�&�;�@j��T6g�2&$�	F)�
a�^�{BsPs�{_���>������� ��~?���f��
i�X�.XT��LV9�	�{�����S���{lkB�(���z��U���.��uOm���BB���~x&�H(Y��J�����ss���%�q�W��L�~ڶ��&չhe���^���[u]cL5���{%��55�ۧ�7�r���s�\Df��R����=+"9>�(F|���.�{5��Ƒ�$�*\�ؖ�1x���6��);�֓V,I�j��v<..|����T.�7#�%h�<�n=���_����Q��UN���|�O~��o���sb(UE���b�"�c4h����hҔ�.qOb������w����F'�F�I��-۝�ŋpo9��^���L� "�f(�Lp"�+���P �9�'�T���)$��C��G;�D��%ԋ	R��6Ct��M����EE2���` ����3�$�D��UyU�C�ܧj\&�c�:ǫNH��<l�ʩ�y��#�����~�;y�/����x�W��p�fsr������+'�6�5I���ا�[��e�?�<�1G��_�dqo��?���å�JC����Ծ�	����#����_	+Sn9z��=q)�u=
:4'��V�.pb J���|k+\����UU��/�b��]��JfRC*١������Ü�az=���͕9f���"��Rm��g��4��>�l�laε?F�����̵��c!�����w儊�`!V*zk�V�lO90��6�������%�Q�{V�7sD}4��}�x���|����ł�+���_}���f�p���rUU� �,LC/�s=jӽ�a.O�����}K����$�c1�(�)�RE�?f�T�����^=RI>�F鿠���M�/�{>�?s��� (����c&�F��
�@^5H�\��IiT+�t�U"�Y�*������
	�&"���Ởj}�=XS�.�.�`c��J(!	<��Ì�� 1;�`��,)����\Nr��}`p�����5�9��	m\����E�ǩ"����p@�%1Bu]�	#��1lkO�pv�cۛ�|�/�{����z����7�{����y�5�U�ӷ�������
��&�w#!��i\��87d=H�l	PS�����:�2]�*H��0X��.��R�����,����=�@T<b��E�S�C�{W0��>x]�B���wx��&X�2���{��t�h*{����ŀ���E����h�Td=��Ӷ툸����5.���$ԁj�]���뚪2����uB4<q�51�2��2��Kn���H!Y���dM�����)�$2م�Sºs����̓*�Q��xB���|��lP�db0e��=���wy	<���Q�*|W�Ӟ^� t&�׉���qJ�T�{��:��+��]��{�d�#��z���rN}��6���H{�s�W��z���X��ͬYS?�-�w�fs�|���r{���]�5���h�%��ǂF�z,�Bgx�*��Lp�vށ�uo�J!dvC��� �K��H�Uk���<�M�K�P�U�40�kV���b騰T��P��S���m�!nˠ����waNA郋c�U,#`ZϦ��i:e���}��1��
+�yGi|�S	q��-_�Ԑˑc��5���Ч �$J�<E@љ�w�4�&�=��B@����d�3.��S�7���pkk��
�/>�M�>���psL��w�|����o����]��}�s[-���uwI�d���1<��Cbf����O���):I|�z&&gN����Xd~��<�S���2���w>�f�;!G�|��kۺ�_^���;�� K��Dƕ��<8u���?�*�L 7aDw3�ͭcXK�<Y�-���F Y)G�"�|���������t�$ ���d�qQ�w.�6\$�_��T�37���N��&�`t:
�K�}_�\��D��"��>m�,���qS��Z���k��V�*^���G�ɟ�0���,d˝o~��|��>�]��%�gT���1Ɛ	�D�>��W^��a:׋�x���1	�b��P'�ݘhiC�����@�0������ё�_00e��U����v.��*���=18W�y:��"eե��̩٦E�8U��Ǥ
���`_)9��{;�Xz��݈Os����*��yw���$x�ԔUM��l���f��p�K˷�7<���r�=?�c�?�s��q��T[���0|p��LѮ+�0��zw���!����5.	�t�����·]M�����+��D���z�b�M���[��L0"4U���t94��������֘�:��YS#b�V��w�H�2;%=	Yx-5Z�G����>"��tO���������~ѹ��=~7% W_*%�O���o��ٹ���N�>��G��ֱX��¾��}N"�q]����׫�^k���~��y���
�ut��g��8g����g�����3����&�(m��pU�����)�p?Y�����r^s��\�w.x����������4gDpy���YZ�a.��31�o�;��Sx��<`k��}?v����Jq���؅��� H��"^|8ǜU>ޓϩ����h~�Fr,쒐@P��b�DT��Ҋz:�4�h"���/�7OȘ�{��{�ł�)/}����ħ����x�g>L�C���
\[�u� z�}�Sv��9�:���e_֟�M:,�&�������w������?k�l���TR`L�h��E���&d�&�������˃ͲFj�T���������QR��?�%�&�כ:ܫ���N�2�O�W�����Mg����9,������'�r�*��ӹ~��\_����YAaC17���5��$}��O�uQ�?Ș�u��ܾ��#ts������g<�<⎜��5����Y���x�~�Ճ�=y����/��P�~�jQ���լ�|Ps+��W��oSC�M��U�Îv�`ZJ�6m7�m����fv`���Nr���%��~#Ќ�}A{��\w�̫Q#9��E@<E�T6%��Fn$���}ȼ�nR�������J��:�I&��x)Bc��]�X=��C/ۄrN�J���;��a�esz�=��3���?��_de9��M��g�[�|�=��B(T� ���\x�}e�Q�?��^Y
���n�$��mp�!��	��kM�E+���Z�7�7Bo����lRi��,,����a>A�����%!���t��2���}j��P���q?���Ra[�2���x��X�s�ɋ��T��WM�;�v�D��Y�,^x%%6�l�W�s_�G�J�z�އ��k]����镶���,�l�������'�+��x;��p�����O}��g8Zm�8�v��2�/>.�Gю��q���uwΏ�ǁe	�gz��>^4��~+ۺ��k�$��k$v좓�t���Ui����H���yN<�n��R:���9/mhFZ�X�~�Y�rh^�����n�"���f){$9��t�S55�w��ŉ�{�}����|�t/=Ks���۟�-��l����'�d�ӱW9�9fgјJ����+���<#�%�����	�r|�2��]~q�#��`%h����鐝-ivD�n��n�l�[\�)Y	�����ِ�D��=�#��*dtw7w^��8���1��c�*����\\����$�DD�}�XK�X�Z�v<ʿӳ{/Du_���e��em���xG�^��L��}kzB�7�������1x�	E�1O���,�ߖ��Ю�����z�G~��<񡟧�nٞ~��_�}��,����I�>�ͼ�'��]�8߾��+s�F��6��c�)R����*�4�)m��ѠKte��L���3��U�T*1J�r�HX'�+�)c�r�T�;w�Ge�tR�K����(	��و�n�?"@542���j	F��vK�B�ڼA����a�̔R�,Ǡ�X�X����,Y.W8u�����|������x�g��Ɗ��w�_����?�HuJ%1q�bX�= �m/�8�����]�������8�Y��0�o�|�s�,�5�> ��?�p{��`a�|^	�C:7Īw�;*�[�tơ����B�Mc��S���o��֙v��N�Q��mJUc�E%Eʚu��S������t�st�����1�?H��g
s}��/� �w������X<W��~�y^���>N��2��g��8���r�ִ�Or�}�_�e��ø�­��%/��"GGX���eiB&�����D��B,��@1�iE����N��z������)�Rx�~7���:O��������V��}�^8ki��[z����<��� iUh�|�SL��i	R�1�loc�q�ݝ��BN9J"LJty*8�)!�
ף�Q�Ϯ!`l\$4cs��gDm�w���T����4|    IDAT�q3�l�+���N� H{e�]�T�e}z���c��ҩǹ�����%�{�|�/�������{?����~飼������!YU gp�]��/�Ka$/B6���ًi��w�r_�a��"�bNz��j�9\��!ܲFez�ĥ�U��������86&X��"->���D�Ẏ�Eob72'���y�b��9D���0�m��g�\��JJ�ĻyE�.�2����Z0]W%bs{u���Q������N��@,|4z��-��������%�+�;=c�$�����a�V�sM89��|���������nr��/��'������b����9+Y�t�n}��p��]�+��$�����q������\s㝮S�}"�F5��n��D�<UC2��c;�l�5]�b�B��7~L����qtY��4&F��E	'L�rm��[��ҽ�Cv:���x�����m�F�>���Y����j�� T�#Fh�kk��X���#���.����`<�+tQ��<��[tU*��1�S�GW*	���]^��NmY�B�U���m[���я��I,�A��r�Ae����+S��k�b����(]r��mϩ8z�AN��5�����-�{�G����_�o��K���?���3�����Q�ͻ/�+��`&�r �1��%S����5��]i��{mĂB���z��b4�KU}ι�����20���<����� 1��z*��ƺ����3I��#5���p������*1�����t=�"��V��C��U ��YF*TM����"9�yx��aL�n����A�(�S����b�Ns�Ho���g2��q[�!�Y�5���#�f#�4~�8>��2���w9�9�]�qnls㞫_��q/��>� �[��N�b� "@ݿ̲]r�3�Xh7k�׎���~K�>J��c���>�я��~��?��{l�}�8�mN�{��j�fCN��X�X�����e;��C��Q���W�dӚ�@/$����.�>�=H�d%�2f:�?������{O'A�g��{�S��l<�fDpELV�W~��6Dzq�*x�z[j}2�.H<��XSŘ1b"/�#8y���u[:	g�rE���o��Ԣ���9M�+P�$�&�"�eTlD���A%��$�M7S5���|�%��δh7��� I6����ݾ�ji��w��?����B�"\$ �HUa�;�;��uO��8��恇��o|�;��x�c���Q�>|���y�l���O�����sn�=�z�b}f qq���������R �5�s�+%wӮι�M��tf��)�6NGb
��!"���"���,���n�ԧ�L��(����V��6l�g�ES#��c��f��p�Oz�+sgh:��o�����b��^Ƽo<W��LM�[���ڍ���M��]u|W�U��G���:�s�_��3d�Нnx�#�n��S�8�w:���}<��[Y5�o?�w>������,�B닯s�9�)�`'��,M�?���	��~8K0������x�0-� ;)~�)��$Lq_�a>�H��Q��N4�GG��s��%���1�lb��8��
D�*`8��r�@�߻*u~���g�9�C��(n�ΰ!�*�E5��uEP�9e���������G���ހ?Xq�u��� +�ylќ�W9����/�o�>�����WO96��e����.<������#��g~����c��=b�������}}N?�:3�Q��wɗ�<[qϼ����WZ;��2��\"Q�xH�_4��Q�(��o��㻽]c��*��~��5�}�4���Y�	%�a���U�����\�򙫔}pQ�w��\��U�����~���9�Kh�c�#�W)1Ws}]���Sc�����ss}ϒ^-����4�u^:��O��?���{���K������/�ܚ�9�둑�[�S���&�O�J��,��L	�.���_�#c�}89��x�dc��s}�r:f˰s�e�0��1���wf�6�W��'9=��_{�0�.o�#����"M���9�\������$�Ka�PnX��}�x�O��#pn��
>��㠩�ڄ:nw|%�F�`$�S`��7���CL/;�����Qy8j*��3n~�����'��g���}��?ã?�k�^>�ik8>�N��ĝ�H�M(e��C8�5�P5y~�L�j��!N���8�S},�+��S���C[���_��=^-�KW�bv73��'XJH�D6NC���Z��u=ׯ_�O��ŵC�J|�{w�}|�����w��!�To_��+����Ua�,1�������(G���{_š;m\4���y/��ϥל�L���1U�fq�c���z���pTs�^q��;x������	/�S���Ϡ''���g=a.����X��7��%���s��d|���ƀi;>��7����t���/��;;ƿ�]������kB�6��U�-�B(�;���(�WD����i2qF~�.Tw�y�)�ɀ�6�J���W.���I�$8Ϸ��p���S{0�\��v���B�E}�ꚤ����f�E�j{To��w�V�n�
�q,��gwXY<�x��>˿.���r?�6���������~�%V���;hs?"�1/:|p9�wa�\�c�nj4eʿsun�v8WcH!̔���h-HS��A��K�Ng{�K������D�	����<䙱
�1� #*X��41v�q�Z1l�p?HJ�SL5��4��ee�`�u���2��Ep>���)l\��c:s�"_�O	W>�0�����Q�y�j��ݡ����ۂH�!�ǿ��,8��mh`�<��-��k�-��?����0K�_�;^��?���7�ƊZ�����Anon���iH<-B�O�<�����8�jF߫Na��u�Vb̜e2��Ic�j]�l�li���#�ᐷ%	�D�5��Ơ�G��@C}��s����c��-U���J�����	;�#I����%���A˃�;HM�#�t�HY�.�1�`P��`�#1�-��+�U�O��U���r~���t~S)�s���B�TU�&�q�e�n��8���.f%t
]����q�3��y�=�(�׸��{9��78�����)�����e"`ƫ�r��Z�I�W˗龍>W�;=k��V������{�?�3�Z�IE8	 t��&�N�2WU��L�ƙ7��8�
����\U�(3��a�5]��cQ7�������3��
Rd�P�u+��� �e����o���i�cZ�"�^E�p!����}�^�`�ƈ���%��7�ZL>ﻳ��U%�{-�60�7�v��B���~�˯xn>�o�͏��������W>ͫ�_����t��༽â1���
/���@=�o2�1���y_���;��PZ���SB�;Pu��YQ���BD����	�:�P�"F��]���� �^@�Gc�o�\CHm0�s4d�Lһ��T;X덼R{1_5P
&�8��yOU٨��9T���>������&��3�Sk�����ǳۃ��\�Ut��CJ�����h�=��%�Eͦ���{��P@XH��札�EЙO%��\òs�՜�9Ձ��,�YO/�Ϩ�����y�5�`��w`�x��#�٣��x̵H]K�y9��i�>�؍L8%�sc�WJUj�R[ꂙ�m'�K���@ ����������{A{�*�!i�H�7���qT1*d�hr�,�.��K�g�s!6�5t��u��:������^��+��)�\T��r����Cq�#�s����U*sƞ{�-<Nd��:�7�u��pIs�ݷF?���U�>���T�4�u����8����}�ߡ��7y�����_�"�=�Z��-۾�Vf^S�J�Q��}W�w�Me_r�^��f����A�P�q�VL�
�N�9K���J�d���kB��>DL��'u�4� `"��L���/Ky�D̃>�Y�O�DU��{�3��$�Ӽ�|�xʕ���|�㞋��|�!_^���
 �c)�����]���o1�r������ҸN�԰9��0O��ؽ�V0����>��J��)K�1��ִ�zJ��o��c��5��?���{�Λ�;������/rʹ`�a��a\���X���y�AH%���M�|������,�T�s
�S�L����0h�xڮτ]$���cLQ�UP����u5���#�Ӽ Să	\�mj�]�y۱0U��q�f0E1D7�(�V�{�)R���J�S)jZ���ڟ#�1��2�{ .�?��\�t�{�	S&��$�Øɍ�_9.�,���E��])r��SFh��r%lZ�{Ւ�~����_�m����6��������o8~��?� ��3��w��>������$�F�����������ŋ�UI짰aLb.<J]hu�v�1` �^=�)}�&�������p'��U��FxLLt�K�Ky]=Du���Ќ&�b���7�Ÿ޺PQ��nH�	X�2��X+tރ5P�u�-B̦�i��z�ӷѕ���)kP�V�^{��C�������U!����@��؊A�w x��B�4(t::�X!G�`a pu�UÂU�n�n���q�Ȍٕ��4�;�%����'�D�CC�q\�t��3��`�ZQ��-���l^�O�߬ꖇ~�X?����<�3?��^}�块0n��m;6��+��s�z��eA$M6DK�$��a�xB���ފ	����=���i7�%��!�P�v��{OS/ú{�h�15�o�k�7!�W�w�>H�F�}`�!���E�`%�!O8"���]Ϩ�N�"�WΫ<���6'���c���E"�.䵎
��Yo���<a����<���w�631N�C��Q3H�R*�6��'MKYr�r?#���r���Or���7I*�5;&��$H$��*�e�6�/�dE��*�#�mbQ���� a�}�$�`L�`L��Tf7�o	;��8S�6O�W쇖�w�k���ݲ���7���]x-�[r�}<s���/��2�}6�|����t�����W�n��Vغ�S����v�8*�t�5{f�f��*��y>���u-q��ĖlE� ��Dla��X��x7�&&�EUp�!4�c�����wx���,��Bwb(m�eAM�P�h1Fp���U�.5�Y}e�5����˨F���Ӑ�Q7�epl�F�{�;,�ѡ&�,��n@�<Ѹ����T�x�L@�RI���1����	�I%Y���j�h&v �;p9��d�wRx����`�YJN�X h�L��,��h@�F &�n�]�<��!�?�k������O���������z�o���e�����U��jj6g��Y:; ��Ũ�!��Hj�uѱd�2HbD$-#&������Z�DN3�uUUh��c&6UE4؞(�s}�0� ���n:�%��wO��l
�4���9FxKsHi�+[d��H*�����A�%�����Z��F�ʎT-vG�8���kc��MIk3��iӒ)���x������13ل L�zO4Y��r��E����j��g/��R��3'���uQ���@�q�1����^pڞ��p|�����`[-x�yϏ���ͣ��>�u�~��|���Ej;E�S�����1*s5�+&�3fpsj{n9�u�Č� 3��3�Π�udx�;kb}l�y�п�aI�������F[���!��XCek:ߓH[�~`�ƽ�k*��-�.2��p��r<1`N�0c�5!%F�c�$|�k�0J�8���%���_� ��O���k��'s�q��h@Dڊ�&� �lD$p@R4 c*'+i� �e�M�T�s�JT� hr�a�O�q��"�G%\���B��bn��w>�{l��7~���9�����}�����6p�>����,�X�|�R���b�<�EȰ܏�� ��S京V+�6F�
��jL���Ce��e�fr�H��1��ЖI֯��[E5)>���8ܣyi��}��� Gy��ȈT;Ho,a���⟁��@���h��%J����HY�֡l{�g8�r&/�<ER�tn%1*cL��dA!"��XG�p�H�H��U(���vb$�S2��u�Ӧ P�Y�_����yi�r[����9�$��+ǹ��[���XXC�r���]�y�)�����_�������֟������Q3D�L����iТ�P�@'Z��'E|Dv�J^�=8��,	}eK8~f4�ao�T�=���xZ�l}�`��Ӻ(�S����_b�����1�#;��F�/�z*�B�h���r�tP���ǅ��~���8ab�3הĆ,�H5���M*����p'���>�$a��l�c܎2F�%1%3(8�T�+�<_)���6�Hh���3��8@�B��}N��/���s}u������'��~�w�u��Η����Q5]�2����9F�>����R�t.;pÚ�$D�s�����{��PD���YH�)�]@����TU���{�z��a�X)��H�4��pц�	uJ[���]�G�L4g�PGX�8��̉Et+e���1��@�t���}��OsL�� ��U�XI�3C���<�b�e��y�3�׋$�g|�D�*jL�(��Ӿ>��=��G�'����}�ߢ�5+��TF�Wny�{�<��_���������c�?��4�}��t~�/0�%��u�,�x_Ϭ�x�cb��??����{��}	��f��0��`�(�l��w<���3\	ހ�kV�����{P#�~X�rCܨ�xq��`Zɉ�ʾ��iu!�ꮺd
H���09WA��%� �17֛��~43���y�[Q��z6r�AU3�Pp�g�A�:BV�����@��",�0�M���b?	[��h�N�v��x׳8?a��/���'>��Oq�����{��y����9Xe�8(�!��K��j��)��O�V%�8ܳJ�!�M��d5I��1x�[[g�/�*���7��E$d�S���$���(�����Ex�hy2L��⤾�J�e=�x�l�ӕZ��$��a-�}�g�s�	���H+��60<�ޙ�%&8�ӧ9G!i�,K�!�\G�1�;�31>��"&a�Q�̧�"R�!:���t��yI���2����3C<S��,���b슃�!��k�q\?Z��ٚ�ۆ���~����}lo��͟s�g��~�7npG,�M��(��\U#��d�x}�Qk��X��4�cN�Q���"������h�C�ݐ$-�1�����B$i�О�I{"��Hwʱ��sO��n7؅�2!a[ym1�B)�dm�N}R��$�n�/��fU\����:�0�Ĕ��$�1�^2�R!8��e��R�ÐuN�4�}y�'���d";aZ(>/i1튠�D<�%�b����&��e�RT������r��)���VG\���տ嫿��jX<����c�g��p�䌓�'��6G�P�h�Urh�QA�݃����K^�bMEB��� &8��,>���Q�:#!�Lb	[�ǉ�.��a���]�"^�F�LFC�wG�,�Fs*��|UW"���?��6���az9�$�}��D�$� �����	�Y���=#ۂhz�؎E��EPu����e-�l;��@ć��hqWzsQ2<�=}��T/Ս�j�+�<S $�49�;�fH'i�˾(`r�����^~ibH�R�U��g_V��W�]��v��c6�J6���j�x�9���?͓��;���o��]����s�g��3��{8�,�ֱ�1�)#��%�g�6�.F&M%i8�E}	׌׼�?Wa��p\�h�.��'�p������9�!�M��{��u�n��uK#����^D�cب��]��<!� c);D����_D��x���� S��$}����9��|����u���@t�$���w�aHm��1ZJۅe2��Jip'ֽy
ɜ1�O�׋d����IkC�$�ko��{_�W�I�W���Bp��i8h!{�d�Ip[|�s|��]S7Bc��_����`��7��<�V�g���>ck�    IDAT/�5F�/-�n�S�����m�I^�s&D3g%�nl�:�S��2�1�K�;����>�˵2x'ٺ?�f`S-Cpg�9�>x 2�딬��2�#��U�!]SU!�}��L��>���.B�sO	��|7�8�i;��,���=Аo{@uG�7ݣ�8�Ü&-�U�Z�%�q�	n�.JeR�r\2�d�!��S��Ma,I����� Wc�,����2�0�!y��rY�A$����a�D���X�Vll��~��x�/�:�?��T�
'������}�y�=��.��>�1��p������0��2�\�qDѼ�����~�C����ٷ�L]Y/=3]��m�Ʃ�:v�mx���a�~ֲ�I�P�!�ee@m ��4s�$�����������`���M7Hdl6z^B]��$JA��_��#��8!��I&,yb�U��ݻ�ys�XZ�kVm�����>2�탇@b��L��d'}"J�hӽl�qg����.R��&�=Y�{�E���6�&g�S����?�מS5X��>����O��?򛬞z?���G0�wy������?�鰦�����8�����]�i�=ڏ،	�àE�Ap��A��,����~�;SE�r�w!>���n�
��ҵ��	��p^�b�kf�2�j�C�'"]Fm]K}	�&��D:39�a��8�W^��8ϯ0t���q�)A�H��S@%�Ü���7&��B�2B���a&lBv�ˆ���WÌ���@
]-�1MK�&�aq���b�\Bb�rJk[M)���1��ރdҚ��Z�}(��^-��Ld�i�}�~a�����g�w9\\g���l�9|����_�(��ѧ�6l��M���ǰ�?Gs|�f��y��k*w��ah��=����9d��`2��v��@�C;��4�}�^I!��i���8	C:-��t-���g�b���=8�:	�͘:�k8�s�����F-J��*�D��Ўb������wo���P��H9�K�ݻ��lԄX�F1V2�mn�γ�m�ǐ��bQ�h*�sTbq8A��m�5���l���m�t��/�eTpbS+!L�B�-Hv���!1ь1X#��% $ӹ�S:����� +a.a�>��W���F*��V���v��xjS�cD6���h�� H�ƙ&�撮3��`+Bc,���W�,V�W��u^}��\��?��#o�`q��O��ݻ��0�@���(D�:M��T⁕����^�Pn� }æ*oi��-A�'W5����zb�f��(�(]��z�a-�[�]�(�N�#5�WʶQ��c����x�be8���9b�l0&��[�^�M��pC��>l9�kV����c�ZX��sf۳4�5�C�P���iX��n���9R��r�*��56͂%5�v�M,����X�JX�p��͊fU��
Z��v=R�cB���`�ϬK�<�p�5�n����	o��mUQu=X����p���s�X�ΖK�s��ؚ�R0-U��9DW5��Z��{*+4�%�z�b�IWs�����~��Vh�s$'�Jue	a2<ueY-WتAհX�jO�<�zU��RA+��9��1l���5�1>h~ꊪW���������h�����+6�F�	�l���uSCݳ\W�n9fA�j��a�t�:V�`t��M��U��Yha�Z=Gt��Ji�%eƻg�\������]R@߰��ط��7���>����~����W^��ѻ�쒍��K��V�OS�s� $�Ӏ1j.��G���ꕘb�[�*��h$%��h��52������$͐,svӕS��.���S�����~XմW1�����RWUp}#]���g�d��x�3�P7uTH
IN����Z��ưXԘ�>&�lUщP�#n�9�l��7���~��l}Ge�֡��"LjX��`��!�w5�+T�����{���,GS�@���ı����Ud���q�d�d�������>16��`��e��KbV��9��Ɖ	W�QY�c�^==u�1Te�,������5̭S���;��C}�1��-�z����x<�	�"<ſ1Ґz��V�/y�+_�?�#�ڻ��#��6n��;��?�w�p7:�e0IyD�+�@���� i/�>�j�jY���;�Y��n��Ε���ؚ�X���Sy���=m�UŁ�<\��D�����,eɲ����j�Z�-���%��hwF�eU{��c�;A]ͪ�0����nt��ܲ�r�����ۭ�ME��8����y8ߞpj�öae`����ᴷ���-���u���W��5V��h�QiCMOc�2xo�\�����!�}��>K���a�*�Kܨ��p`�ҩam�"��>�u-'�1�lg�[0��hI'k��n����%�kײ�k{�v�ϕ�o��5�m@�yǶ�,�q�(��5��5� V,�3H︹�u�]�SYZ��{�m,�k�����Y�#���Vjx�∗��4昅Z �5h���[�Z�����F�|vJG�rQ��5��S/�^��]��dK}t���ܵ��-���im�����^a��4��ǫ�]��]r}���d�[��L�8"/")�^���o`���y����W>��_���Ӹ�3����.��v��U�����x!$�
�[)	4�.$�s4ĩ �z76����}�:���ޒ�%�BP�x�w��˵��a��ϟ��"���$-UX��=\<ܸ[70.�YJ�)��4�r����x!Ŝ���ʚ7�ʘ�o�&7>�f.�H�Ub�Lpw*��U���}��.'����
��hc�u0d�V�F����{�`��	i�+{ONY���!�T��f�́3�!R�x�s-�kH�P[�áV,���gk�]�w����r�_E�-�m�����/5�(�v��L4'!T�"��B�T�">������;�I�ӗ��cO���O��wZ��2�}�#�đ��e&�D^#�~�(��0�c��%��oў�bũּb8x��x�mo�t�@*۠F�^�l���D������w��q=�ز>?�z�kܹ�u�x�[X_���4,���9��1�[��s�Vv��n8��*/~�<�[���۫9x���������5���7�������z�5��q�{���醍}y�}lzS��9�����1�ca�;��՛���78p-5-�Y�eQPcYw-���=B�p��94H��ځW,��pG��+�׾w�#A����:D{N��m96K���2Jמ�/<����c���L�7K�4R��^a�;|#��CNձm[����1g��;Os�6,�����؃���y}����b���Ab3�E}���ZT��k���RK�,t����+7_B���uH��.N8ඩ�����Mc-��;���t�7ի��b���P�H�"EY��%Q��m�������4�'�A# @�!H�Hw�N�A���nKjI�LK�hJ4%��H�S��*�����g�C>�s����`��](T���=��q��_k��2��(u̦�бbl M!�5��
�X@o���fbbY��D�$����c3IiI%(�$�BoP��*!���2�s"�+j�p	&pZ�&��,L�:�fv�O;K]{�^����*7wn�,��2���:���H���R�%�>�p�]��~W�SzW|��@� kC��20�� �i
AESKλk�]�ѷ��4S��3g� �Y1efl���_{��V�O�J�Q�ڍ�0�х��ߌ|m������u�H0��Z&��2�cϼ�5�h��0up�K)�y����x��w�kv�Έk��D��;�VS+v�w����;M`Ή_#��pԮ����~JD��=����=��`�>Ό��o�� �$*�x��������ϱUt{K\w�A6Μ�tC�1u]S��%��Qĸ�P���)�T�N�ŷ��f[!�.h~�{�a�`�����I��Ïk���z�cu֯�ΛgW��R!Z�`����m�?�'K\޸"��K�N��7���?��=�(y�a��HMhc#������[_�2k��DW:QJm�(�>�N�Q��!"bc|H���cp��TU�t:	~W[1�\����'(��{�i����laT�z�M�E���I�ׯ���CF��s��*���>>�qY��N�[�5N�FȄ�F_�fo�&� �C��/���kF����H�KR��v�i�M�\��͂̀����x����f�����ӿʡ� ���Ғ����'R1�ڌ)�x��o|����c�V���i��S.����x�/|���E
�1>���$J��ls���;�#_}�Ū���!�~������:�:�K��DR	�f�Y �C���&}v���#��?���G��E�d$bv72�C���^d⸜�sR�ڢ*��$�x����.;O~�~�}��܀��u��3���C�"��q1"����0�*��|���c���;2)�Up�g����k��=�+g�w{l�����o��*v6�p�[��z[a�2NȽ���C|�4.��n�	'��<�hs�Z��L�q)5�'Q��[���a��p��^�3���������Dƈ���{��Μ���7̎񬜀Y�5�*xw�j�+%�{�l�k���4�+��P�K��$�g?Ecjه��Zh���勣u�{�ՊfJ��O�fQ��bߕ~7�A�B�����gS�*�N��8����x�Q��|�3��Z�UN|�2�z&�����$��*�)�R��"
�]1�*6R�Q�#8���^��|6��+"2����pPW�`��ą�
z�H]�,Im}��q�����p��+vg�@���X��N�,���ef�d���1xy[{}�ͮ��$�;8YS����x��?�yW�5^'�
Q�A&
�C�D��� ׽�!�Q�JJ~�%u�\��ja��?p=khƅ%�%F�ʠ��jHE�(�X��-�R:)���>����#�n8Fv�0�Ê����\�Hz䱥s"������6�{�Dy朤�I��ㆇ��]���1y^��
c!�
g�=���^���2'�p�+_`��ߥgs�q�.��#l�g���m�R4�m�	�ep��[Np�#�p� >�D2y�	����Ș�X�Z�;��'0x�����g>MH1�UI�S��"ѩ���ٿ��nEEem��!�8'�"8�?4Ǹ����3��WC�$ê�[o���c<#�BJMY�(�㰯�N�}N��E֎�]A�����w��r��c;l����Ǹ���7&�K��U%���0�`L�򉣼�ɸ��UTT��!�"K���P-�ʭ�7}���>�wd�^Rk�cޢ���|��D�ʋ������kꆦ~���=�װ�g����w{��qJ)k��q��?�}FyNT�)�}
<�� t� �Q$J�A��N�-�m{>7�y�}������:^@YW�ŸHN��{,�	��ڴ�QM����प�-�5�=��'��v,��&�t��&��Ț�<��̃��!��0I�k�{)v�om$�.׶��zw[pgLedP�B�]����֢����F��Ch3;�{��6 ,t��6����n�{%_DS�Ux�-�}�VTZG�C�D �i}�Ak���!�8|���0��Ek7��_I�q�Қ8�"�����	r!)�y�F��n���K�:���[�*A�5�nn"FC�͑� 
�/�*�a9�I�l�<m���3�c�37J��B�&�nq��;6�t����6X�&�sF�
h��	��,��.�(2�vDEA�i��C.JֶΓF��D�vl*�T�Ex�7�s�����o}��� Q�Z�2E]�II'r�D`,H�}�H����`�F�2��u����=�o�QU���{�-�(����NY�՞�j_���&!���������|��8a�6I�"�',�c���Lmu��p�}��y�9���̓�fD�xr��p�Ϧ������f���H������Z��w9��{P��2Z�O0u>F�sh,��K���*��9p��M�y#�C.��W�a���c��{��}��%�O?H�6Q¡]�9A�0��K���gy��Q��ɛ?�=	���ۗ�"���(��gkjk�Jb�b0�FF[Fr�(��MEu�2�zIԃ�B�ս��}s�я�0����5�|�*�ͺ`^8��D�d�n���~�����M߯���VY��s��؇>�(��p��IT���S�WQ1`���s
��X����0m�u4��'.��❵��so��W�̞ɻ-����B��VlW;8�Ȥ#��$�^�mk��B��E�5�ub��8��
B�]���*GK��!5R*L��N%�J⥢vm��m�Ԡ����W�k������i��FnL�E���^4��Z�p?!?=+����*���7G�>����AŅ�PbZ��
�%X����f}+�'ӈii:gޚ&[Ρۜr�8����e�߽1������b��(왠�����o�����vMJ�𔻆q-�������mNm��Ds�B�e[��UDl����B��	���$>����Q+M�����qz��@���yh��<?���ꁋ�x���n���m�y�\^~��~zx�ҽ�s�(�|�-�5tY0N�Al��F�zG��	��͆),��,Y�k�V�Dc�
aj��ﳝ�_Tx�!9�t���V�l��MOl�f�A�TM]r_��jd%(rO^Y�QD�笾�"��U���e
+Cuĥ����C�<�!t*x��ˬ�?��3*o)��C[��W_��VQ�A	u���:�	�4�	����x�'�'ۋ��2���G�� 9L��]�C��3o�.��.6x��Op���sHjb�+��	TW!㄂�$��B��Hm�C ��$ғJ�Sv���ء��=�C*A1�d畿"�=ZƌG�Xﭾ�'�/�6(E��Xs�����aEG�]%,�S_=OU�$cL�4��{⨇�}Lw�[`���k-Ϭ���|�]F��C�|����d��b<B��Q� �R�(Eu��ŧ��7�M^�c��1�ǲ�A�2d�I����+��5�X��سv�u��ŷX}�5E�ˈ��}��>��t����d[��f8"��Qol��.�2	�����g�m�^{�*��e�<��?�Q��<c3�WW�6Gŀ/)7s�A�C�=�	�a�(��~�����L���ݫP�M�5�d�@ʾ6�:����	���ڔH<����&MK��p�2��JBL��Y$���K,���U/pZ㥦�zX�0x�����U�DTXQ�S�I�RN�����!��M�e����d/Կk��w���Z��Y�D��Ѿm:�Ӭ.����ڹz�{I�I��+ŵȺ�~&,8���Fз�R��V�����~��｟5L2�l�4�h>T`ӳ�o�h���]�����y�P�I�o6�j3f𼈦ߝD���R�k�Z<�$9)�ux�I���>R�ǎ��������_��_�w`a��{���k/<q�ܱ���{�]��9�z����l^��^yyGhb�{�7���b�<8��,�j8&�R�^Ba,*NpڳQm�	EڅI�/���a�RzNhR���YT%�Gz�qV�&s�h��`����券~�7��CV�z�e�B���(�(�#7q�g#�-�,]�܁��1~���8��r���8�/?G�{T2�h^�qV0*+"�饚r��|���wYs{�ko�'����ĒHX9�o|��ͷ���ͩ�c,�m��@J���u��p��'x�����Aݍ)�C�1QY"���}������}��s�!�l����y:�K*��&�C�;pm�]��[r�6`40�5�DJ�S�Y:�.�~����d|�,㲠O����X/-Go���?��GU���8<��3�K��دr���b��Ć��广����`�A�6*�:x�?�҇?Ψ,�z�xj�ށ�������2�%k�<�O|�z����F8�8��)*O�;���V�ޤ�p��6��-SD	��[O��,ʄj�<�=�8��*c_')R�#7p��3w�9��    IDAT-X��n��ӏ~��j�+O~�V���>�'��o������\|���iw����D�����ЯS�s��>�ￗ�m���EV^}��z��a�Q!�V��sl����]��Rn��Y{:2�+�q5VY"初A�I*guM�B)�Xz
�g�n�6��F�Jj�P�!#�N��`�l0O�밝&ꤨ,	n�|D}�2ó�^��6�� �Fh PR�\(5�1�UlӴ��:�V��Kr���	����/.lo��j���(�n�9x$�3�yϖ���$��"�("M������0��}�P�F���*Ip}�х��@�2!����s�җ���2��X���
�
�x:A�'�O`I��+�Dh�)|���e�����t>�8��2��:�A{i�GޓE�p�E��!�^��`��dR�f��ܑ	���4�jiH�&6���A�(1Px�vo�?y�w�k�7��_z��g�]�Ж����y�{��_��9�/��<�u���%����ya�C�Do`\&FE�oH\[�FH� ���^ �.8�{�ڔG����D�����B��
hɅ&�Ա$qc�vh�b���[p��)�f;>�+=���(��k�x��t������(>�xK1ԁl���j�,�����1���kɒ�l�+(����c�I����.��=����Ě8��b�x��Iq��BTھ��61�\�x�9�`��M1rH���#�R8�0~���U�r@�Y��bl��l���-�Pq��~����u+��{P{�m��HK*��K�p�)��7x-�UD�;F�iɐ�؉Dr��:Cl��D��r����07�D24�H"��2Z�6oT�����c�,�����Y:�a(��ݎ��ȑ�<��װO=����U�XFf�x�5^��݋���c����Q�c�������E7�Hd�܏ @�1��̛��Wx-�츈����Л�p+��&Gň��P�Ⲓ�+t���&h�r��O���>Oq�:CK�KL/"�5��^&�2��__�:ra4�SG8�����:��ċ�n����O��W��W��әgd3�0GiA�D�>N8�鿇\:D968x�T�'�+��
10L2��S_�,)O[@e��@m�$j&���s��Y%@	5P�Ld�,6
е4T0��c�0�-$N�H)IRK�Dƞ"�� 9q��c�n�W�Rh��J��cI�Cm���
g���Z�m���D�C�`�YW��B�T�h���8��EC�>5P��r��t!���pg��O���97�G� �O�
���n}H����˓ �I��p^Zk��B�Y7�h
��8נ��f�y��28�I���2Ӥ������&AY��5�����.���	1j��럇k��م���sOk���:k=XQ����Qds�����,���r}o�DK�ǿ*r5�]6@S��M,�v\dS���5�*J�뚾����a^1\:�y�,=��׿���/�.��>p���7���:u���i��2���.�Ҋ��
�E��>��UÄ�;C��Y��l����h���͘M���>�w:���}� �exJ�q�RE9۱���%��8_C��1�5�(��*!���	E"�Y�Jx�zהzĎ��)\(�G�N@-��ak�����F��%㔠rM���T�B���MrX�F)�k�k����S!�'I"��C,KV�o����&Ne�DR��Qi(\�V(� ��x�<���!��k���QH��2�jKiǁ�I;�XP��->�S��Qe*_R8��%��6�^;�ҥ����Bj�h@�:�4"W�&W|�ʥ�,8K�&X��8�$Aynn����p�Gn;���E��UP���T:�p���C�+~�:Q��}'�O�H��l�1�h���/p�gоd!є�+!����^�!~�r�%^���3>�c�$,ت7���ƫ�нp��c'1�&� m��\D����/g�����/�VW���+c"�I�Bxr$g~�#��/0�����tek�>�j�;�a�Y��d���w�.�u��6������i��5h)ɄB��J�V�Qw'����9v׽���2��ҁ�I+�(�Έ�(�W�*Bw�ˊ;N�`�r��g~����T;ۘ|��F�*�R555ƙ@>$RJb����'�@���4�cԘ)^4nM��>c�V%���P�.���g?cy��9h]ծ���� �q+�ӝ	#�M6�>}���o���^~wP^{�O�w�@�禼ح@>��b�k����w�y���3ʡZ�!p47V;�V�����bB�[��Z;��H#p:�zd|dt�g>�ٝ<����ls�|�w^���88��'�ٮ�R�+OS����>���Jc���������v�l�P15w����;��8�>���-V`���#+Rt���NPUa�rS��A�kЊb��v�,����K]j���
�G{��@E�-�IL��S�*K���נ������iD�IZ��K�1"�@G8�B]
g��!tH����	9�Ьc�k�B���)A]���U5��X+QB�ʊJ�8'������	JR�{��eC
��!������1���&ւ�[���i��-t�s�<���S�Z"�#��)�%�HQ;(�B�y�\�]�9�::�>U�J5�F:�T0Ϋ��e.%��O���������"0VP��\���[ly��o�s�C�|�]t���A�WT���/x���%����^SJ23�/�K��2f�C���r���FY`F���i��:K4Ũ��3��'�-e�#L���}��g����
�F��$I3Jla�D�	k#�w�T%h����:1qՊZfO��6�7�k���ٽ������0{އ��=�=EY2?�ǌ��ܐf��s�&n�;?��ݏ�@GԖ�J���I/U�����P )0o(n�������P����Ս��yš��s��g�y�������%�=�?~�= ���	ʉ��Z^*�����3�wءH?%���Y����ݲrw0�ޙ�[S7����6�R+���I�����؏��7ȫ������o�o�}�]�;i���3S��ɳ<���y�3�P®���%�g;;���]���jj�ZZk��i�_��Mn��^5�J�W�V����u�Y�����_��Ǣ�'����7h���/>�ԗ����痾v�I�z�p$�.���F%]�Nǹ(&�3s4+�w�kyD#����^�]��u}���(S��;��.h��$�Z��qc���A� <���q'�w`	!#��Exo�h�1y��)Q�ol�\J,3t�֠�ǚc=^(��H�R��Ho���?�r�<�uh��P����0���1&�F�OjԶƋո3�s!�Ӂ��<���@���e�qΰ�l�yTةKMF/�4��T� ИXQ����u!��ܒT���������Hg�EbqJ3�5��Ա
T˽���l��}I�ua���ْ���,um��멊-����yK�<�THd�Pc˂�˂�/��|,-3�_��9j�p;ی�#�	�I�o��;��GJ���wp���		���٤�a\�E��j�Q�uO`G�s�d�{�����UE�r�MD�4�8Al��-R7�@4O�-ua�H���*��d�q�����øNL_D�5Cj���U��N���vϼ��v��ݛ�vM{��<�9���&�Qd���PBS�)ä�ܽq��f�����r������&����5G�����0������ϭ^8�*�d7}ⳬ>�4W��s˒|���!����M�΀T�0+��*4�8� �B���~��\য়��
-u��f�'�;��s&�ج���ό��Ϛ��@��zv�g�m��x���}��,�Y=��(!�M_���޵�E��mA/v[����g�L4��k0|G)��x�0��`����8��>���m��g��/����� ���]����gs�Oax���a4�v&�"dTx��;�m�	�)`�E�]�q�����I��eEl�I��KO�
UaM�1��� ��8f����c�D�S
_C�!�Z)��p�蟺����o!�b�D����G�y�n"�s1�&$u�t�(Q�IaJFC���C,#�PTΒ�Px�����(5�;���U=9d�u-��vA�IS��0����v!%��Lx���/#��4�1�����t�]�NF���T�1O:�Q����g��c�˗Ht�lP1��Җ���C'�v�25�8&��T���{2��;dYOb�q7C��;�ֹ&.FQ��xgɲ�K�m��DQ���x�stJ�]�B�:�R�B��UW��8�������\9�㍯�#rL'M�G]�!�H��VH�pnH/��E\e$�>ȡO|���e|5$�^�����^��%��^��EĚ�ڣ{	�h��vd�yVkϰ�����ȣ�:|����oS��:��D���2~s|�%�{�w�����O�ҙ�K�n�H� ��ȗ������3�Bt��z��_�h����O�����S�S�o�����������rgtSqDV#�9Ҍ��,�69��y?);u���݆;���g��U&H�>s���-ں:'�o/����%��>�?�l��771l[��2�:�v�5{�nu�r��������'Z8{�����fj���Z5��R�-8�H&��5�V3�{:Ғ�~�d��neÅr)���|�	p��kv�[+T⨬%
*Eq�-������]��5��Shw��o|����_~��-���C7�&��&�ϾET���m�ۄ}i��g��
�IQ���B�0���B���g����ۭ*��q���ct�E�� d��5^�֒��xz�o$,P�%I"P��kF��b8d`,y�I���GV�kI.-uO�[y�gƗ��Qc]�1�k��0փ�����-<I��(B�	~���zh��D)�0!��;��O�;Z׏RD�F��a�)"�e	P���ﳘ�������:M�����B�qs�������
]�xы����W������EɆˉ�<���(�>C1��,�y��?Wvj�Ń\w�.z�%�('K"��#���
/b����C�a��B��2����ZT��4�K��b���xL��EDUz�H�1l����s�bH9�$����7���~��.s7��"W_z���e��P��4�f]L=�����r�N8��ǹ����u=�:'���ݯ��7���9O�#(�%�(��Ұ������X+,��9���9|�#�� �&���l=�4��K��&��l��z�&kM�λ���T�m����v��j15�hҐ\ңH���an��_E>���.$����r�҄��d}���Ο�=�x��� [?2�����{���E��)|D+EgϤIܙ�e6&mj�5qC�us�?fR�)���n��G��{�I)h?k�O��� �%��G���~����a��ҳ�Z�g�t��}�V��T�}}�3����T�6���I��:�M͞��z���x����Z&����_��ƑjrO����0���P�3��Q���|v˃�tߗ�)���?���k��]>6�4���_}������������W���ZrhHY�U3es�{���\ٌ�P��gK;�9F/��o`��Xi�ӘHgx�Gw������,-3o��c��V��G^�1�),i*B���t��5z'��SvjG�-Bi��$�кg��`��j��!=�0'�c�^�Sz�P!��[�U��6��9���=�dQ����x�����I�A���Y��Y$�nbX\��*���;���Yl���*����KK1�Ȣ����K.�1��P� �5&/0u���UʲCZ��I 9��G���r��>�\�c8ޡ�=Dl���OFY
��'��8)��@Z�/U�o)|^�P��Ұ�T+\G����>Xe�-ҭ-��K���6��;\����8~�}���A����<*������*�i/�Q�T�^w��Q��q����,w��/]�L�_�����3Oq��_Ü;�@�P]QF��%i�DIY��q�S�T��Y��C���ǘ?p�am��o=Ε'������<i������}����"��f�����gsأ{����I��R]��7}�Q�O�����d����?�����J����a_N�����{�Px� C[���4��������!=��Z�bZ=�5z�qy;3�{�a�C4��{]#{��:5X]k47���L���1�UK�낛aVF[�;��u�K�xS.�Y~7|>[;{V�ٻX�����T)\H�l��[�b��3A[ja��-��=�w��~:�B7RN�&���uj7��~6� �����Y�7�L������ãk^����������o�\������N?���5d~!(IM?�Z��s��nv3OZH��M��6+��ܧm�tP�^2T�r�ހ�`��[Kt�vn��_��{��1��C!���f��>� ��2ok��*g����D4�O2��t#I\��r�5���Jjj��PW/�/�����"bOeJ�%�#b�%*
E��ň��b{�^8�u�c�,u]���5��M�tzX�0u�s�uDK*#A(�.p��v`�F	��Zg���s��_�w��	�զR�J�	Ѹb[<��e��-6�/���k��1#�#|m{�YZ$���S�!�9:�uQ ����N}�ȃ��\�X\��ͧY}�UD1��;(��c���x��g�J�D	�IJ�SY��Q�)d�p%Bd(k��a��Y{�u�:�B1�:{�}���n�
����ddQ��<���'������Qɼ�0�1,���oRc�^:@%1ۣm6��������K�a3��V�p0��y�_e�ų]\@����1*�7"b�puNg!acT���}��,}��~�B:��e�>�4���'ī��&	�C>*���2�j���������b�O��F��8'�`yc�x�i�=�Q��'�����/����я�����z����lQ���z��o�8�U��5��N��ک���nJ�lyԩ�4��w�71#�f��k�M���\��ȵ����-��V)a"ӌ��f@׵��fpX�5T�5��R�-�I�5q�>����.����Hi*g0��GH���kZ�M�>E����d�l�� �P�Ϛp��P�^8�JD�Xbl� .�Q
τܺ���D �Lh[k݇Xt��BXGVzw�b��;^;y����;-ԟV����������D�����'o�|mĠb1�Q�*��X"�x�"��Ƀ��cm(�j��i�`~@���mn�Cy�=y��֢&m��Z��� BR�(���
I�$��|�1�N��qX%�]I��PY���ۺę�>�����@���d^0:º!���������sxS"�N�������.NH��@%)�s�d �mR_�T���*�ga~�$������@^s��Ӽt�y�F��I��!I�G9�]�5[$��ʠ��.GzO.2�0�$���A��J\���k6�}�\�����\���C�^���%��4B�R��q<���B2��dkc��A�$[�zI�j�z���R�T!S��1^[|
�Ze���7W��E.��<K�;"��(};,�D-0:fю�-
�U=�ј�#(E�r)5�m�A�Im���0z�/ImF������v�,�e�/����Av8{���:���;ԑ���H*�a]D>V��z��>��|�n�(f�M�7���7x�L�\�ʷ�;a.��1�5�9�����Sγ�?��G?���}��G�9IU��	.}��a�z�O�S�xH�<&v"��=H%&��{]�{�Ť�;�w3��ɇ8�aH�&�w��GA�e;l-�ħ>�����I�����m�?�����?�����#��K���ӵ9 jCE��"�U��^�Z+^H�$�ڄ�+���u�*d�D�FK@8T�v�	.�^�0���hr*��q������UѸ]m� ?�kk��k�/�� ��9�B�d`tRP[A�z�B�X[�g;��Z�i���mΟ�lv�\�sh�n���)�a%� �V� L	�F�p���U�)���H��f�}nۗY��Z�]������ dl�(�    IDAT	DM���<e��t���-���&�p�����wΜ?�/��Bv�f.\z�2%lV���M��݀T@U���s��q��W�8c�J�ܟ��=���{���-�h�����C.Ɛ�V�c�#�1�Pĕ#
���l�s�����7������i\� D�Ě���FY��R�xo�bM�DaC9�s����t -N�5%U=&r@)�F	�l��1Z	Mm,��"��
�JP�5��&����Q�cz�Pz��(�QQ����Oe�87t"��3vʊ�:z���ի��
΁��(߶|�Ra�A��H+bl`�Z��%N�P�R�F��A��M���t�=~kL6��s�O��S�rjp����$Io��xH?��>��O���S��Rrk�ӖaY���J�[E	[���غDT��bЉA�3.$���D�)W�u�1�Qwҥ9��q1BǊL��!���J��êd-�r��p��?� �6C���������_G^�H�k�RG�I_����.����e�u�m���C�p�c?�YX 3�Snr��g�x�Y�+c�J�
��	��5�H)������c��'��qBG	޺#!p:N�>7�u����?�t���/���n��_�헾���N���.��2��y|Y`#HT06�1X��E�hH�0��NeU++�u5O���Qq�%V��~�i��J����?3�@���ֆ��& 1��� �i�0!�Y�oc��[G�쳿�Z��>D\+�m"'����S	C&<��D�����d�Ƅ�����Rre�f�vM���S�_����]�@5�X��9�=t���$xoז����7׭�G����<J%eS�$�P�O��,�����B4�G���2/���"h�3a,���a��}�_K)0��,HϒsD�,Q�(a>I)kC^ٺ|���7x��_c��š8�(
6\�w�'I�T#|��s�/���69֕X[bMEm��҈@K8�b���D#���K�;7�z3o>N�E9E�Jh_������*(F�rH�0�DD�$R$�#\�����`$Zh��"FTW�L3�
(RT��)ǂr�iÜ��IK_V��Q3H#z���Qt��!�I��D
�(B��"�8"��,�פJ`�JJ�$c�����?����*����{�'˲�����{ofV��U����<�@X�(��$H�p�V(�Ѓ�:���)��� ;l:a���IE�4� @=��檬��t���9��{3�Ѐ1pGdU�ΰ�>k��Z�B�>'�قi�1.�[}x@�c�(��s�-��ak4"9�q���L�h� ���3�s�����P��9~:����w��Rmm2�aIbp,J=����:�l�N�;1Vgy�/�'>�>�OQ�,n~��o~��>�G�o���f�b"�aXVl�)v`�p0���������*͹Ӡ���>�'�ē���_d�u��7e��j�d4ap��p�C=���ˑ�w����!*K�x�1Y��D�9s����sW��_��"��[?�!"z�Ƶ>:y����y��HN�f��֪�׽�7jrQД�����2IU�d��q�Ǻ�ۻ�;~����`��׌q9� f�δ�B�걘�~\hk~cTD�B8Ǵa���nW/p=&q\��o=Y1�oyZ���\�W1F�	Jq���sg8q�En>}�y�!�bqEy�:�stc�����fu���r���.-��k��z��y��ߺ�ȍcW�4y�/����>������ȣl�� ��&Ng�&��Y�V7^�@�1"�,��SK[��H̺A�ʱ���F��e.u��7qs�%v�t����P[�z-��nf[�nL�ٝ�@Y�dN3�18Q�g>o��o�lN3�P�m2QI�1��kL��@�H�P�j(p3��ll�:E���A�0s�P
��=C�P�#�(����d#L�h��B�F�8 hA�P�%���8�s����-s@�X�QS��a�$�&®�!�� �I�`f���d ���=�<�դ�Uӭ���Q���Mīgow�kWw���ޭ���}��@ʬ6ݐ��TpE��1ej(R¥@"76�m���G����Q+��g���c��lp���};���N�8q��_b�C��3��S�����~�����!R�aC#-��*�U��Mٳ������ϛ?�_s{� �;TE`�ɯq��>N��������/W���4�5`�69`����(���/b8�,rf���c_��O}���K�)�����sbʝ"�Xc#$t�����)�&v�r�uC§�M9!5i.y��	�>�:�=��"��^���Ƈ���w�����{��>�!4S�	P7q�^F�\��^4��"��[���_de�A���x�t�?>\�C"w2 �Y�}�AY9�bd��L�n��P{��Gc"�e-��E����0��X��zLq?�X��E��Y�p#���P�ΕT�����ð��a��q��9�l�*����<۝�o��rH�u����O�f��ӯz�o��+�?�ȣ/<@�}
?�Ŧ�9;~�E(���Z�wq�L�%)�1O>��6!��3���]W����O�>�����c{P�'���g�����0��0��y��>�3�K_�"����J1E~�c"�^$+��	�j�XJ됶�fJ��/�(�F�뚦�����Fe�{]03����#�H��=^������u�F�L��k���Q�E� o :�|�^���#
��'K��ԓL�u���0�H��4wc��Hʔ)��
��5�j�)`��$,^{�'���/]�054��^��_`8:��<p������������N�������c��B��f"z�[�������]Fi�a�a_K���x�#����]�3#��9��t�roN�yo���1z�[)f�u�"��[�}�ٸ�2%�a�S\�|�~�9��+�&�fʼ�RĄ��i��Ʌ����#��6���6W��&�|�/�>�<�!��2�{
�j���p;L`:e�m�7-�;u���A��L<eI:�����7���>���/q�ڤlQO�fbq!`b``�:��	;FƮ�����ݸ��t��k|��q�gK��'�M��鷾��r��?���)�{��`�O��/�/^|�^=&�M�hH�갮<����w$�s!�����so��,b�ʲ��r��=�酣�q�+�f �܍�H�k[�n,��m3bBS��qݤX+���;�3_����h��
���#�Gb�6���:DT���k���'N�g��34��$�YZFK���I��h�A���~B5Ǻu8�^���y�|�2~ۻ���ט��f��Y'�R_}�2�EH��#�U�%ѳ�������!�n�u�]b�r�
�;m�nXkIQ�Ƒ���ւ�M�2�ؚቂ�����>�<T2z���M6_�F��q`��d�bʲ�,*�"�b�ÉA���R����di�� <Oe�����l��Q���؛�*���x�[o�co�*���8�a��L�k
������	�-6)N]���N:��M�J!JC"F���u�{�[�N�.�]���0q��_1/Y�/�^�ۆ��uI���R�B.y�~z����QPF�R;W��dTV�n>��OͰ�q�]�@<}���S\|���8��gnq0S�HڻN��"�>�M���6��ޯs�����ÚL$�9�
|�x���s�bNr5?�63L}H���h\|����2�6�KO�D���ࣧ�x����{��8�"q~���V�mþ��zy��w�<o��s����c�mq�ɧx�Ͽ���+Xw�m�:��0��D݄�N�x�,78�mFox~�#����	2�r�{O������.'��xqFj�������35�Dhj|�qDa�?;�L��g^N\�N�n��WUQ�> �Ór���e��7���~BC�ѿ6g��?��b��%anr΍�)l�r��Y$w#��w�{��tBv軚�eE���?��]��kk�0.8ꤾ�!��g�Q�F��	�Rn�p*�I\ѹɥ��~r�x��1����U������/~��Nwm''RV��>6Xg�U��t���M�xnJ�:��DX�r7�q�/���\�Σ_��W���| �r�U�P�N<�V�'<N����S�_���%Μ��jk�5b"�V�c�q�G��Ү��0�ƴ���G���k��U������:�,E��(;��u4)�S������g��op)Լ��=^���&����_�\g�>���f�H��4s|�	�S!`L�{\G��a�f��8�	%ab"�q߇~����n&���i�"���� ���m����K𿣗/Ѩg>�2<3d4���i�����7���.�y����/a�
h	�D�֞Ѹ������?�v)4)cA�mt0+1�e��8z,�HȈ��_|�4$��fFJg�h�rɘ�Jy�d��K���?��~��x?��!��#�f�g��O��)�s��>�i^}����no1|�kx��{c��R�B�#Tۜ{�u�a$��������T�]4����Ë'a�<l�����[O�cvs1�̌� g��^�����-��un?�u6�����~�x��|���g��P#�a���I��}���n����V-ÊI3fs�p��/0���p�?g^�f�m����c�}�C���&:���x୿ �����L��$�P�e���~�34���8��Zn�)�;����^.�r��.����jPDL[Y�m�.\x�շ�����~��&|���[����x��.���X �iI��Q���js�Z��8�[�xT�[C�G����\꘻����y5e���v��퓘�4sO�Z�A_w���1f�������භm�^�W]gZM������!"I�N�g��fED� ?9dv0Ξ&K�h3�����	�n%�o�UR�NѯS����E�@��3<@���V?��Oye��v�]�c)���0&A�5��W��֕�"#Ar2�S�;�i�䨫���o+���M��$0��w������P)Xd)av���s�Y�5/}�	����[~��z�;��l�j���s��e�<Ʀ�~%`LKKi�B�)E���W!y|6��"�'8��7r�=`�US��g20��	��Q]|���܀i
�pHAI����NΦ�Aɬt̊��y�a��2O��b(�PK <���4/�٧��>K1�6���,���Qѥ��YՃa���l�D"HB�!i�H����QZ%b	M�$�I�O�(��$��Ol�5� z��	��3ݿI��g(�.�KL�-�����a������ބ��
��M��&en��}n�k<���p%a6�ɿ��cx�����#���|�k8�����)����4"���:�ť/��~��y��!ψ�8u�w��>� ;�):��s6OX^#�g���ҰI	�mo�*����S|���w�iN��^�������f��-��9BI�9y�g.��j�0	3<#`R��c���O|�8�pj�uOѯ����A������9�����\	�Ery��`�����O��G����������'���?d�>�]�@�.pa!康da����1�]>^Z{}�(�����.�V�uq�ŵ��%��G��؜��F#6O�"�d������e�lJ��$�X0JM%�&��R"��B����>��l.H4�e.�cG��2'PJ�p�:�9���H�,	���W
��k'��[�v}��zRH��V�-�ZX1 .�=Իˉ��8g�i���e:��3<��.��'4�a����x���������2�sbj(jGr%14�|E���N��dr����4(F))EQc�{���w����K%��Pf�'�3���O������2x�)f������f��[@�=���׿��=��{/���wq��/s2��-�}��l_0z�ܼr�Y�)L�9�mqlT�9��3"��G����k��k�۽Ω���9M9��Q���F8��xLQmS׎{Ű��rjtI�����ܶ3�������ov��$­=�7��g��S�?�4g'���i0��TXL��4b-�Ѭ��d��h۩QI#�Fli	�������()yv��ő��Zʀ-/ljd�ҷx�3s�;l��}��8�Q38��-+N���n�Oxƌy�/~��*�9�1m��V�d¹�M��0�����'����(Ԅ
�3��a��q�8N�)g^�(�Ҳ�5Z��-�E����or�����>[�n�O�K�N��5g)�4�{7np6*��1���0!fdP�$j���
�3�rl�#q��F*�@�5�møQ�D����i4�y`�T'Z����b�3��]��,����&/t�]�	�
B��(Z�$�Y�e��Uٰn8�������о�BN�b�Mh����������*�~Lc�����Տ����5�j{9H��[�\Z�$�����;����ζ���2��d:Q9v���M.����hsh�ҋA[�YL��BTO�jk�����I0�� 5�C�>��l��$G
Mn�e*��CC5��/�45��:$@C"Q��vK��'|�[������u���{����`��%9���8}+����,'X��JY*��G���e���BaX������mmRG4�9�b˲���Ab��ۦ�rm���N�껵����'����#G��������P&vwo���ϱ;�3���ᗾ�;<dӕ�:��ߪ̤F)���d���{�&ݾ�y�ӟ!^y��gOp��_`�[�y����cs<f�`b�u�e�9��D%�"�P:K1o(Iؐ8|�)����r�[�1�ڠ�3gFp���3}�;��uLc�1��4���ͯq���3��1l@b�U.�L��`�3B����>���x�SFs�&'
�j��>7��B
	��,��69ve�W�2m�ln}���_��f�|<��g?���yr���'$e���F�]�������Y^���p�w���n�0��q��&\����y�9���x����[�}��%4�ٻt�g>�G�?��ݢ>s��
q�`o��c_�֭����p�k^˹ӧ%�s�V8Um0�|����_���2�y�=g��=����_}��g}�3�8����z� ]�x��H҆�#'��^��ߒ�7�x�n_����9SL��-�f��AN��L��?�Z�O��(�m]���'���5,0*�">2�����Lj*W�ʂ����9�p��}�_w��7Ə�>s\��yN�:}�}l�<��8��d�j���,�:�.H�KN]蚮!L�'Y������FZ�y̹�a�6lK������x��s��m�DcLKa�ן�7I�����d<�}�,�|.�4]Ag�*b������w�����k\��l�G����c��z<�(��Q��TU5�}�����#�G��JMڟ�;��xá�U8n��N�j�v���Owl��>M5� ��mw��X1X�0	J#Ęulǭdo����!��0��Apέ��;J�U�ެ@cV���!�#��N��b2=d������5úa�(>f�
C� ��#�����U^��? ibxv���)w�0��c>�-f���҄�(>6�M�u�ACH��E
���ʂX���9���W��/�}⛘�c:�ghqI%�w�{;Ր�I�(�M�y������-.'r�*$FH7\.Q3�)��[���M���Is��J�i��ѧ�C�˔���S�$8�e�|��<��3P{��!�KC*�I͆TD�9�	&*�d�䫟�矢ϙO�(��"geo9�N��o��\}��_@�#���X*k8��ev�Y�z�V����@��9[(�ܾ}����f��2��\$pN��D�I�3~�Yd����a�j�b�(7�"���ع���+0&�	��Q$N@��R���߽���ѽJWPMw�����T}���_�8��8���T
m�Q�� � �}v���w���L����N��q����O'x�����Wn�}wx=��8'���&1KP�;E��]�3f�/�F#UI!Q�~F�2��e��R-,�`r���M�jf��w�%��Rѫf�(Y5���    IDAT����+w��̎���!�EY�28�[��:�]'�h�]۶�v���4g[��AW���R_W�]���7�h�2�p��V$��������1��c:%�������Uw_���{\\�5ؐ�4M��G���wC���6�pEٛ�%}W����,�$ �
��ba�^W���{6�y��.l�
6�0��L�G!� ��9�j ZD,�hT�[Z�B�B`�p��Hb�:�~�8w�b�!��-R='�,�׭��KU�L���bҰd�RJ��z�ޜJPjh
\Q�B$�����آ" ����k*�ICjn��!&��Q��"!�t��kF�-_��1�@�he�EUK�Σ�'?�h�f�׭��$�l�9V�(!MT&�Z�P1�!aK��F���n<�e�u��>��Y3���� ��w���7�u`8RX��t
m8n�p�O�h�bn]M��Ԑ'KK2����\~gK�)P�ך�f�a�h���st8]lS�֨���t���]�p6���p��H�c f�04��Ec�h��-��;��K/p����ۊ]T?��9ԭ�&L�@"���a��K����	�%|̃~pBBC�t6���HUr���zh��\��W�fF�iF��x���h���$�2�K���\-��p�/��HZY���G2�7t�s�!9oL��#FZ��C�u���k�4��l�����2-Hj�:�C/}E�f�ѷ�
�Z�*�"�r�H�(<��=�1^(�E��~w���}F���.!��F-�.�����{�������h����ݛ�/>|�����y���UD�ɓ�ܙ-
F#j��0���e�%/w��wP�ݾ����ܳq�M6����J�1*C��DT
B��N1Q�Iu���}�XGe�a:��8�� @�SY�j.����	1�l�w᝔uCeI���F�cs�*u��F���Y���;(I�Ш�V',Mm	�P��#�k�C�1IEYRb>��;��MC��gƹ�11�|cH-���saeI����1�@�lf�Zr��i�{�Wŀ�'��1!yl��� Ua>nh�b#�g�:z0�qQ�U�(�#QbX��b�X�8'���hy4�2����J�k0D��d��y&&+Ή*�@�a�,�*W�Ϊ���1Dt��s�6��B�·V�%�H���%a�c��XN�<bZ�+	!���A|�-�0)b��S�7�����r]���7V>pH�u�yB�����gSUA)|\�*�s���uo����-�����4�ُ�l@i��ٲ��J��Q]:"Җd��x�N�s�w��N��<y��
��+��h����젮��S܇�������tH��[�~�X]�E�Z]YKsj�,��I�/�����rcݹ��tV2ˉ����Y.`�y���jh�(<�-�����?���Y�?p%~���eN=��w?�/��&�(���ic�1�b��7�k�e��â
�=����z�!����+�~�9��rP�!�Ф��i�P�!�@�x
g0UI='f�B�MdPLE�z��4p�
�����O#b�����k�&bj�
4�tĔ���)�B¬�)"$��i&\�D���Ԑ<Z�$q��6e{O�FS�	s�gV�"&C�$R�PRUhTB5X2L�dŝ��'����O�3�&bmr$��R��e2��Äx�@������T(Y�
,�(u���\Ye�"x���a�H�BR���.��k��D�-@"6��3	�*��46�Y�M �JS`.*�G�d,!hC�u3gP�&�40�>��kLĔ����msU�*�X31�f�`
�B���
�qV���&GT#B�5lr�/_�QW"�"��h��Ǯ!�Ǎ����Q�Qs��h�)S��I����Χ!RX�5�$4T��Nk�m���G�ٍ�kۑ��s���ި�)iEL�Dmݛ�ém2�B���AP�ļu�  ��J^�J[� �]������'܂y�x�����}ȡm��(��j�h�:�c�BLkհ
�{�w�/����,(v�ovQ����L�w"+�,�^��'�f<+Կ�|Yw>�F�ݾ���K�V����Ԇ�O!��.f�9&)�q�m&n��s���^Q�ie���歵�RľG�q��N����R��d*@H��-J��4�z���*ےɀ҈�:j��X3ĕ��sj�)�g@��=Dɐ^��hgrj˰@���Iur.��ր������Q��ZdnZ�i���Ȑ&V[�R���CR���)n�-��B�x��$���cH�u���Xr 5>���UqY�+"cta`��ZF�
wQ�i�����Q		)��aTU���מ"���ihNҘ���kc�e��la1�����F����	)B�hH���:�8�1��S�D��W��̢�x�ĀG��b��(���F^ D����04�{���X�b
�N�h��L�NP�ih(���[H�{B�>%H)���ز�4S��W��?�Gr~~j.}�)R��|Y�$PWV����}���su籭��E�*��7���+�;����+��ж�m��Kj��O��^8�-�^�&ۣʥEx��<tQ�-L/��� 3��^�w��ލe(N������UY��BU��]�T<�2�u���!V#�������<�p�;7�r{Y�rt�����RK��F5m�r�v�H8�o<����:*�C��@����.�����;T�gK�g�w���xx_�DQ���?��|�-s*��xWf3�g�&y��0Z|�U�}�`XƎ��}^��Y����v���A
�[{�M�	u=gdGDͽJW �e�MR�pܞ��P��$�hľ�G�>6r�<���3\Y�>�Ĉ)@}Z�JP��@�XtF3�l�HE"����::��Oi�V���º�D=�1N�p���s&�	Δl�6B^'W!*�(D�-pN��s C����	m�&���'�+{<����A I$�H�
���an�SN��̥FS�>�n�4tX���fP�&�a#Xh�y3�(
6F#b��fư��M��`�`���el��(3ߠ�8W�B��V�'f�)!E¬�J)J�ڣbp��)˘p������DR�2�ZnˆT���b���R�efrY�%-�ēY�
�i�TE&XjR��H�u��Q��W�w#�RU�M��D�l��kޛ`�}_���[�H~�8%9p�r��&;;o���S�нqg|��kNl���n:�d٭.���
0;��"WS�ў>Jd"��*��<O��eǞ�:֕|�z.eO_i�1��>����U�&�,�-0�U�2���ة�]@�`�r�����$]vaJ�m�8cQcH1���D�}⚤i��IJ0��ӊ�t�B&�i''������[�c>Fl��:{r�ߔ"�DD
Dr�}NK$p6wpKm�����1,J���{�RB$.>��(�3fD�Էq�_���<�����ql�e��x�r6N��&�7��s���l��ͱ�D��#�� ,kwI{i����+̛�i��P���n����E;�v�;�*���m�$�ɒ�*�6ֶ{-�|B1��i"q����EΜ}� "U�	��o<_�$��g%�T��4i��,�5fd ��]"?��3������ mZk���!��L�2����_���߃)�xJW"�}.}���=�U�Y�4`��zƼ<���]<=T�������)Jn'�R\XSGr,:�U��ڇ�%�Rf:ˢ�a��"@�<�@i
�Y�J|��=�:nϔ�[[���&��wѭ��i<�,[')Kǰ��ao��7`L�&ŹANJ�])�A�ŧ�\��׀� ���ܸC��D���uB���Q��fnd��BTC��y��Ts��GeT ��460k�P����Un�UP�D;#|�1���H�1�el,�(
�Qʘ1���e)���6l�y��q�[��{��� 
��}�`l��H����;8Jːg����{���\���!��
�O1���ߎ����Ƈ\�Dl�̪U����Y&�e��"�J�\o�|&���hXP�y�n���%⣂���QST��ź��p�|�|ܔ�-�Ut�L����5e�c���ڐC2 m�H�٢"٨5Tq�$��k�G/��"DM��U�K�|��i�bH)a�=���� ��ZA��0�'����묟�<,���2՜Q��.��`�ya2��wq{n���[ά��|߆�r���ឿ���Mu��o���$?����jj��4���,��-v/_&̦T)R�cN�u�5�7Hg��R�t���e��d&T�	b�DT[س�_,���4��FM�A��
B��r�KFb:��}�x������E��q�������g��@\��Z����5e�l���JY:�������{�۸��8��Z�!��^�:S?!��j����r���=W�7�eAU��|��6���XG��#ƮdhQ�n=DYd�D�R�i�4��Fq�2��N�v�t�`}�k{���u�m��c��8T5C�k��eB>FFܖH�q�AT	�WU�19����y�&�{]����,�^�cL�We*����y�?�ۯy0g�&5��|��w��w�1Pؠ ֺ�
���T��D��)�޽�?�{�GMy[O�ko����<}4�ò���& �|2g{c���?����b�{�?����?��ƀZVy����{�Dv�/�mwS���gŬєrC��#+�$���˶@������K�_�~�ر�^�=}
�G���)%4��Ik�^BB�@
z�zF{w����R+(��	u�����?��P��9J����e���E��C�Df&�.���-|�mǳ�kHH�O�7�ݺ͍��5C?2o�?9���#�?���Ƞp��p�;��"2�cD[v�eN��x�Eh���v�?����i7~'���9�s��a}�t�����0Yj��AQL��cZ�C����U�Pnm2�k&S�6O������]E\�7�+���5+d�(��h+��>E�8��`����A�s�s�f���Y(�3�Ulq||�o��f��9w^������W��`�P@[��z�������F�F��7¢��<D����'�K$�)B��uC=k�M�i��X��+s�aZr�\K��ݧ�Q���3kY$_gl_���F�佒Ĵ]������-9�B�in~$X2mr6r�}`�
����ќ>�ޠ$�9Cu߽�Sg�EA����޹M��m�
��5���;n=W��ů����#�4o�1{��V�:rbTq�{�8{�����x���8}*|l|����� �J�w���^�Ik��6�2�����}n���Gs��a����C�1������N[�;�!��d}�C=
��"М�nDPY&ӭ
�la�׻x���5kq1	}���}�������댆�;G獚%Z bZ�9�����a�bw�=�@�C�p���>��}���������Q�?��]�c��q���%;�?��u}�)��]�
�0�5Hh��bK�`�%�IG�h����F^�TX�`=�f��v��
,�G7����[��%Ze��0�"	�2�<�A�i�̳��0۶rl��Ɲ����g���1�#Er�y/u@kJ	;�	Ed;0�%�>��\n�8㶸=5��ݲ9�9��a1�%�,�-��ۺ��'�4M[t|9Α{X{o���5E���w	�w��B���F�>'P��)���@��WB��1Bݐ#-RӢG�gIDr�k��Y�r�pڭ���Ψ/2,�P
W�� ��/�I���a�����ҳ��u]��>FT�96��l��v�P��Jtr�sDg����Dڪ��%������#�+����/�ݥ��=�!���QG��w�p㫟�W���c��ql��_]����A&���j-��yQ�ea��U��ms+�Hr��IA�d<cH��){�=�(Z��=�_�IߝGo����bǍ��%��	�-3`j�Esy�t�k���s�0ǘ�2�7����ȥb�N]��Z��N�g�,�2�`����y}�͊�ůw������nd2A	��DRj'؂8�Y(��\����Co�����7�{�������,�׾�,;_�
'^z���L�P�Ν`{I�	%�.�.+�~eD���b�.Yj���uY��+���]}^��m�����Ʉ9�¶js�Д�8�FL�3؛�綴�-
#9�Z�c'���?�H,�mL��-[cG�0P�L94mR\.�1NIMn��bHuf-KQ0��,KF)Q��5i�}`ot!��OW�t��q����|{�����{d��Ҝ�$�h�Q���c�ň���|�+q'Nbc�v�mU��i��oC/!#���v��c�R]ܯj�֓fedZ� ��ܴkIJ�rФ����&#�u�յ�Nz���S���;,�Ո���4����!a:�0Gbȟ! ��tɧ��GX4�Z���hN���F�F�E �Ξ:�ϡ��s����
K�<֜�t��K�z����o<��3�I����;�����kz�eHx�T��j��q(G�M��b� �C��֧y�rɚ�8hϹt�R����[��
`�	4���^�Ӓᨬ�#�<L�y%H�P��po��xb����
�'8	%�&�h[�ߝx�\ޤ�RpZmK��6c=X}�gP�Rae�v�ם%J{.Ŵ0����О��$fE���}�vԠ�)�ш��2�
�_{��O�1����RU�ZD~�e�܏8B�i�9��7��6n|��g����5"Đ2u��ԧ�*zRfw�J�ގ.���g&�}������[�����W��;X3E�y�ˇ��6�$%����E ckqEAH�lx��	�/�dr�S�H1��3�I��LVd�&��[�
h&��n���|�SQ�u͆�$�`8s�L��P7�&&ꦦ	'�Z��q�nz/uHٲ��e��XƎn�w|Z�X��Ϝ��em�hM��������0z���8w�89`.��$��s�W�ˠ����6��`�E�_Qp���=�fi��9=#�{��n�P7�z8�9�e�M���9����QU,&�"4���=="m��甪��QT#��dh�n ��z��\�ݗ2�ܕ����q��/�ꑻ��X1�~���oh �"�*#vX0�5�7O39�e�k��w����~����~�����?�<=��w;/>I}�&#hY����F��t��fi���ޝ�X(���eI�&'�J�	ֶ�ĝ��##��G���9zc%<����X�u�����"]&(��2d~�iA�{������M��'?�	�R�vlkһ��w� v)`�V_����ߨ�(�v�!��w���>���e6�,h��]L�.�����5��"l$��j���9��w�����?�y��z�/E�ٗ��?ܘ�����{W���_}��gW���Mf/=φ��[O�ㅅ�9�>CF	�Ѷ.�ͷ�N� Ԟ2�^3F�'�mEW-��GM��IBAN�\]�e�UC��2���S�D�4�BVC��X�q�f�Q�qdmc�����2�R�o�k�,;��(���X650}�[\-n���4BFS�O=����h6V�Y�IK�t'!�2_,?�����P�#�4�;�bȥ����g)#wX�u�\in��!FH�Q��w�����g��8k�UIq�:">�|��"x��BZo��ѻ��y^q$��M7
밽�k9��-	f�װ���
�H�{:1-dCH�@�!JA���W�ɥ�B��{��9n�)1-�x�g'X���߻�Uiz[�̝���T�y�8<&D��QC=�f��h{�_[��ﳧΝ���zfwsj�-�I$KTLEp$%B�Ȁ(F (P�8����{�XF %@�`æl���H���f���Û�tΩ�=���wթs�}-Ŋ
��N眪ڵ�^k}�w}W��C�Ϛ���Pݫ��_�!"�����ݿ��CG��J�$�&H�!W!��t�ؐ#���ؤ������ⶍ�T�1��7��q>�>�b\Ǜ�v�Sζ��N���k�O�sh]*�
�p��+�_�#2UʬF�g>x鼓���&�����x�rX    IDAT�b�<��}�y`�����Q��H5�L03�>\�0�MN��I��$&#Y�S�JR�7[�tA�`qw���v����מ���?q���m�����{��ι/�5���{�s���y���m^���xO��������:���0����ɖ�D�	�r��(�U�0ARSF��9e� �6��'QSe�b�R1&�P��1_��A,�*DAL��his�jw� un����+�[q�>�Ѧ<�YN�\�'*e%��|ۭ:����Sz/H�w�2F�%	{z�׿�e��濢�kvU����Y�qqݳ�7W�PJ����Lw��|M�ѐ��1�<;�n�i��0>��|�6jJ�hb1��,��x�&+�)c����TMdyx���%��J	�)�Ύ�H�$HFf��s�c!nHz��69PU�o�2�oK�"�")F�9CxTcN���	�HD+�٠5�Q�i��RUn5�Y�o�3-A|��5UV4��@�Bjj�ɪ�u��.O����ṛ�yd>���Q�Q�'��tӸ�Nkj*Dt��8k�+������[���o��� ���Zn��?�G��?���_��k�"'K���U�j6sJ��L)�&	�q��C�Q��I�LQ�l5ka+�,L���r���Rx\zg�?v=z����m��5�~��Dh52�s��(�Qv-��F��	$l��2�o2��@J1�$rĬʄQ	c�B�����&�dŨ�]�ǜ�B4)΄"4%�O��T�Q~麦g%~�H(P�UY&Ԙ�T��mP:����x/��)Pt������g��Ou���,�饥1WQ�����|�k��cҍ9���|z��0t��,��o|}��_�
�9z��n]�����퀲-*t�n ���@���W���M�i�qD��2.v��{�����I�D�y�TE�gS�q�3�"w��by!I�֢%�L$Yϩ��v���2��Ԓ��V���h��hS�y����
���5I%����]b������z�	�H�.�1;	Q	RTDjLo�c��ː4+�q��3\�E���ΐ��<������x�{���a �-G8�9��~Am����:���7�#�X,������J2J!����u&�$1���Z��&�QA%��P7	Z"�Z�> �Ak�u��֠�E��$��}����ۜ�C�}���m��	_�x��N�&��Kv�|�A��(�(�&��[SS#6#V�
�JkE'�%K�b5u��C
�oS5(�@�re,V-�ɳT�HU�f�SUTE]/0VL@���Ƅp"�]CRx�>i��+������j|�XհV��si4q8E�
S9ZS!VѯN�>kߓ����&�CO%̈́es���v�u��B$
Y&�lx�*i��1���gd�'����db���c "9������2$��8�(���÷_������s�w������������������y㥯�OX������TzSU�A;����D�DA�8��,%lTU�7�T��l�s1G�ر[a��F
��*�����!r�PVŔ�TKJx��Mq>3qN�r+ڂ���I�%k�hZEr!�a"������.�㔍>{sO��%b�t�/1��Ӟ_}�>���M��*R��(���H1���� H�<�1U���%*�P�wN���?w���t�0G���\{�u{�>��}:�EQ��(��;�ս����]���z�/~����ۯ����*�}�iCǥKX�.I�N��Z��~��w���oga�4�"؎N7�-,��0x3'�Є��&�C�X؈�5Zvw#'��b�k0�{�rUQEM@ʽ������`[BLT��UZ�C�]��@�z�:�FE���k<R)- �I���e�����ݖ��!�����1Ri��B���cT�`׎��@�Ղ�(N��T�f;)0t��X۰��ǥ@W����E�+����t} ���!iM�mFU$=v�J8Zt�J��ZE��K�����5�$!6K}�1JpN��
�^�l�E���Z�2x�hv*����&|�a�c!5��%d�*z8&ƈ3�+��T�z���gC����·�I4��`�-i�B�L	�9��;���5������º'&��,�.��O�:�	X�(�r올��DT���RE?1L�IB$f�C�0�Y��1M��KC��mK=��Mki���G9�A�J'Ŕ6��nXӶ1F�a���&�����cZyd����{��w�q�&�;A�3��,�U����x����p����}���_W������7�~���u�������'�n }�B�c��\It�4���5V�@�f��.�S
�k�q���������m�?{�x9��I���a�h~~m�=�����a'8}\�Ș�+�G|���W��.��� ˌ	��N�l�s]ޔ:���م�O�,<���q�D/N%�K��(k�ÚI�#:�r�V~�$��;�N$�}���U����������g�x��O8����߬��Kw��u��oN�n�����o��W_�C�.�D����n~���
��un[�ѓ<����[�|>Vgg�y�yy��7EV&������3�K�P�.�h(�[��~�Sv	f�5�W���Ի����k�P*�����X�=K�3'غ[q�G]d�L)}S�rG�\r����AgɟU?��t����P�����,V���Q�ϼ#�ce�J1�5��)O+&v*AU�^7��� �h-Y@Eh\�Q�n��t�����@���$���w��`��c�Vd�80�i����;>��A�(�k*�%��c�i`�9��]n�ȐZU��j8lk:���xpH��fĔHKO���{���#;u!�ƞ��%(O������������DPˈ޻����zRJXW���%a��ڠjAiO0, �1�^/�]C��S1���v��=֘���ɍf|dG)jrI�U��w� ��:��UOҖ�*z�`�wr>����X'ϲ�h��m��qڟP7�̀r7BI�Ka���q,[V����4Z�]��}�c��>o}Ok��i͍<�(sb��V��s��7�����^4��E��L��;�U�;���tz�O���S�������7HGKl�)�1��&������>�T��9w�����^���0���6��y�y��)�W#Aoc���UA�TA��9@f*zނ���>��h���=?^�"��1_�CiS�RvH.�!���$JW�� ϝR[�J6����HibS�s3C#*���C�T)�H��^O)c���d̿�ޙ�&2A�6�;��7߀o�p��5���s�y��.~��v�=[�ſpU���y��_����}6�D�~҇�/�8z㙗��3��ηxP"t��^��=K<Y�<�ӄ �$0��'l�r�F~��Pۿq���{�6�y��3���]��D0�U���4�&b��*��mz�7ۧx�Os����V��_c+�v��"��w���Ǆ| 9j�چ�N�n�e9m����O��>L�,�Ւ�r����^���?�NZ*D]��������7��S���NX�=����Yv�@ rǵ�|���>��5�Z��w��]��~�}�"�����Gy�ß�z�!�)� !Pk�DX��np���w?�ò>^!�%�[op��os.W*��&u=J)�J1X��MY���=�8W|�^@��l��5�n���#8��}�������Dv��4�$�8�4'WD?�!.����6�!�9'ި��O����$ڣ#N��j��-�_x��R;�3
֜���� �?�΃��]�EZ|�[���Ap�PUBw|��k���U;�g�9��Q����Ԗ�`��0,.�C��t^�"�c�M�b���DE ��]����*�[�B[c�o�>܂������!1�Y=�Z���x}�[q�D��()��JY�7M�h������cMݖRM�hKH���<�����T�E��u��{ܿ&$>�ߣbe1�	�Bղ��Hi�p��?�ś��>��z6��������R7�+o���+�����y�׫�7����g��+�>�j-%Dɶ�j�IU��������pt�Q%oUŁ��$`Ή���J*sB�%�c�s΃�X�s� ϯ3��Xg<&�H)*�[o�pLF:Ȝ7[�)�D�a��K���1`è�<�?���q8=)䞺Z���ez#߿<(6@��H�ӑ1ݐ˲T�$2�7�lV@1�s/._�D��Ǳ!��e��hrc�--{NV'��H��Ex�G��@��C��'�~�ٻ�;��nղ69RJCǲ;���u�;�	wnsyX�X�^����?:$uP	�Ez��/��[�~ףW'Rr52>r+��m���(���K6�9��Z2>ϕ1�4���V��K˱j�y�)��Gy��?ϕ��˩�,�M�22�Z��.x�	�-��heIX���&}�*O|�<��_�3°:�>}����������ߧ]�1ڠuC�<����_�w9�*�Ԯb'�r��n��
��anJ���S?����ٟ"�������w<����?z�.��^;���ӿ��\z�Gr�WhJc���!��T�Fb�������?"}k9��p�U�7h�HңTh:�X���8����O��aq�AN�=��k*lJtC���ZN�x�ן�׾����
�wG,*�`+�b������/�G\Z��ʩ�2Q2B�耭j�{�i���$��>G���]]�[��a��ʕ�e�zz}�#����������b�"C��%�F[R�"CB��ۯr����n���o�z�(�zX�A�w�����D;���|�o�M���gI�c�^2��ᇘ7Sg���_{�?���'��۴Iѧ@�@���V�"T�x�ӟ���>�8�*zT��B�=��u^�����⁋��.n��Ԗ�oۖ��jl���0�Ҧ�u�m�Wrf}�	J&}�-h�L�r������H��N�mE7t�(�USs�����|�=��o������_����>����P��߽ټ����������'�?��?֝����9~��,�z�/1,�R�Q2�<!�M3)�@U����s��ض�,�%�]�����=�tL�n��G��(�0����3N�h������6��NG�G?#�� �yϕ�@�2���IR�}3�,�CP����r�WFe��Qd#����-W?�ޫs$s㜬l�Y�#��%qL	h6�q�EǦk�D`�����x�yĘ�G�`�U�V+R���m���}�l�@=�-��}�`�b��4)xb�!wV\2{z���[^{���6�{,q�����8�Yv�b���zd�r.I���v$�G�ܓoq�����Y#��r�g�"S�S����0p��>�q����Ņ_bq�"��N�mU=D��´C�]ͨ�g�$��"C�G�.��n��bo�z��D�p}��^&V;���� jE��n��=!RGp:��^i��+��U�<=��]�-Ƿ�X���F�7���1���ʒj��As�П&����5�4�
V���x�k���8x�w}�a�������vL�v��EZN���'�d�]�`.]�oi��a�n�|��&����������k�����왜�_!<��c\|�	����*�emj*	V~��-.�:n���:��k�΂$
�jRR�̓<��'���Op�Ϡ�H�O1�*�[g#�B$��{�'�B�����~�ݓ�$m�2P9E��O��O�|��'�ͅ'ރ�|��Xu�"�&��,1z���޳��j�&�?Z1)��e�j�D,���|���%�ʢb�D�k ���~��x�����|����r���\�m&W	lBM�ѹ����ENOO999�2���@)UHaې�|����iMO��r��>����4:������gO/`iX�v�b����W��O^�֏�j�����>�k����~���1�籼k����ɴZ=�>��ٓ��/��ߵ��W���w9z�%:�R$j�j5�6`�Q�ޢ�AHw�M_�,?ځ1����-�:��j��l���4�j����P$S�ϋ�a���5Ϯ1��m��T.p���w ��|�gIdrH(7**H��u3 c��8"h�'��Ű��"
��TB�X��o'��f0����P�%�5�s'$M5��@a
K�D��>�4�	R�L5�W�Qj���1U��}��O]D��q���2���t�]eQ�C�A�v�VLn���,���^ᜡnx�9]���!��� Z1����co�i2��g����l~/r�6���<����7�g,�=�QH��+�1�o'�<������O}�Ԭ� 1qɵ�Zac�u��5��>�@�霯jv4���_Q�Y4�ݶ:!p�z�Y:1y����(B�Я��@��ҭ�Ǻ��W��ĈE��%��$��b=at�g5)�S���i��`H!�k����ʩ����
�!��;�S� \����c�x�+��?<�?��[��x�����#?��<� k7ob��^�h��u��5��@��$�9�z?W���|����[���,t�V=m�q�*��TzD[\j4!�`:B���ɿ[ߡZӐ8�wİ~�a���s����-7�naRG�0,��4�E��2GYq�,v0.|�c<�<w����i�"�k�����ǣ��i����Q�w����^���6�0b��v	�tDE���㩏~����_}��Z�s.��QP^��p�P�H*f�7�T��*U\z�x�����У�prD<9FV}1"�PK�[ETFIN{��k�f�0�Iڴ�Ós}�|f�g��XC>+�>�ƕ��cX���$��%�ma��Nw���~��%���������8����u�=�Uu���}���2��%��orx�du��OVK�W������OOٓ���8h*��JV%[�@��JJrZ���k��D�}�1J�<�����K��KÞɔ�\[��n�?��m���A�?��9k�m�*9�5VP(��A�1��#1޻�o�ob#[+��4Զn"��L0��M'LŞ��An�=�1�w6�t��F�vv�сP:3�sz ;/Y�S��9����q�~�?�m�+m�F=���Q>��%g�"��X�#�I�ԭH��F�"���� �Aeb�Y,�Q8]FH�8!�!�1�cH�R#k�F��������^�s��:���7z����G�&~s�P$/�Z)$)|��͂t�2?�O<�臼�M��Kn���;oA}����w�ikN5D����z�j�u��gV��ۼy�m�,O:v����(Q:�R�G7T\P{X*��k	���&�t�c�Bz�u�+�ĺ����*R{�K
�:����TҲ
�$�KT+�hT�q��[�rw�zg�����}n�Sg�!q�>���{|�g����t'�I(�2,�y����{��p�o�pq�Ry�,WHߓ�*D��]v��}�^�������������u�ђ*�8z�G���\:�t)����Z*�i"4��KO��I�:��5CwJ|���k�XKoq����G8��U��ǧ�6E�Mv%�p�
k����"�ʥuIs���?�Y�����wn�O;vm�����>��~򳤽]^�u�������a�D�g٭p�zX�]vv���	N%X�ّ��r��)��$�g@3`�����,R;5ڃ��O�{���3p����&�|u�>��,wYJ)�t�GGG�q�eV��C��gS822�g�ks�6�次��������d���CU��@J���X�Y�ĉ(�M����+���?���˸��_F\�`/SM[[N��\G��ݒ�:f}�#&!u�5�>Ѵ��Vc�RJQIpؒ+�A蘇��qV�@Jt;6{RJM�;����(uWk�Q��n�`TM��|���"C{�Z��7%B�φ��Q�v�Խ��*�@\�)?�!d�$O,�UV����6�IV�d�UmJ�&p�%��c����B��$T&7�Ц�L�H"�mT�92�'��h*��$b��k$d�nI�Ky|P�����#X(��G�#g�r��k�#�63��3hhb�,��U��U��M�	儔<���5$	i|�*e'h.��H&\��rmmdD*Z4���ʊ��.pN�v    IDAT�TrY��4r��x{ږ��}͛�2H�_�'jIÌ�$3ORJbI�?ź���#��|��~��X��1u]㗚Z����7x�w�̭�~���ta��O���^z���t��s{�����7o2�:b�X$q�����B��e����m������bҳk*����XKM�,���h��
�j�`1��x�F�9�qƱ�
�r���{���-�|�~韢˩_q��'x��?�_�"�4ʲ�V�ء�����p9�$�Q���nh16辧m�.�g"o>�%~���GV=Q*}�}<��_D?�A�rE
�9%��=~�c?�W��\?�Ǝ�H���?�/�]��.�����'�K���c�Uo}�wY�їX����:���6�	mױ�G�y�s��`|�T�Zѿ�?~�+���k�Mͣ�������`�`� Cϥ��|�����I���ܼ��~�Iv��pg}Ⱦ�B����:׾��i�w�֑��K���}ܣ��Y��څ!��t"����B����0P����4������_���C��x��;�������O�M��քe��	^��F'�9����Q)@
��!>pr|�bg���s�'�ڶ�o��g�n���3�!�
0�ͳFk���
�FD7%[A�t�T�(-���f�#�L���o�4�@Wu� �0�q��c;V|$&�X��
QBY� �/Qs'�q��褚���)�Q�<�9tU��,����J^R.e�`U�V��"}��DT�s�@��\&���@5���&���|��uQ�M*sj�G ��V�
��r�H�r�j��g��1�����F�lT7��ǭ��1/$�闊��K�a؂K���~`�����"��f��Xѥ�~~N��
�,>����-
7��M�-ͼ$ #@ܿp�B�+m�9��G;��\�%E�H�bܘs���3�٭|R>�Mfg܆�d�/y( ��n����n�2!�2?�z�S��V��&�BT&Ed��R�-u]3C�Я�����|��?�΋?�z�5�!wbR*��T�F��Ի��R�"��8�L�(����p0��h2*RUFi$�ҋZc���I��S<)���Ο�	$(����2��.mZ�m)���E�CL�������7�C�7��o~���H��3�KW$���ƚ�Z��Z[a�&s=��d�*�!�s�:/?�]���%��i~p�7�k�*����Б����q�ؽ}�| =G�<���	XSM�[�\����֍������'�^�q�O�6T�A��`�^f��R��wD�h�fu�o|�Ox�k_���1�v���ÞT�s�'>LG�J�Bb�`�~���%��6->�Wz�薪1�8S��[o��s�D�y�6��]�J���4O<
�`k�R��i�^�hPP*o�����k�Gvh�� G���ы����Q1p�к�=�~���]y���2�FU��6�B�gL�	cTFQl�!sɝ����aoo�F��:�M�b�������{^08��z��h��h5�H"ab.��J!�(
��a�f@�B�X��/bH�"(��Ȉg�����C��z����E��'�1�!y��)�9�,�UDJ�_�9�i<տţ����l�Y*豺g�tDlRJHx�1�E2t?��B�!Rff8�ߺ0�0I6u�
��]P���M%v4<�YԘ �#V��5��[�H0�u����L���������DR�`�l�)�)W��1wV�x�[0�L �\�Q�S2�$���\�|���cy6}�K�de�j�ȷ���P|�旕���[���;�(O*w�gx/C>?�:>��nCVw�U�����
?yװ����{��z�t|Ⱦ��J��B��M��!�Ecꊝ�ss[��Q��(��R 52����`�<��(k�^>2(�Pv���\��;@"���Y���Z�Җ��>ׂ[�ڲ��t�Lc��o�^��u�&���8��fQ�P���MvZ��>���G�t��SWC��}�E����ܺ�7^|�'���ڊ�N�hQ�UC�X`��)���N����Z�,%�UZ�@Z\j�X͢s��}�)P�
���K.4��}��~��'\T��$���~��o����8K�#�0�Ȣ��^8�OYV7`������w	����D	�"��i�%�@8`y�����p8!�����Vo^�JS��E���Q��N����Tq��G\n�b+H�����{���'��/���n�vQS�
�Ae�mI�E�Hh�P$bt]��*��8�X�����v��`�6���W�6{��<��Q�V @���k� �����9�)(pɧ�����n"m��:5f���9"�8�� =`%���0�������Kv�Fw���p�6�>:�YIu��R�4I�Vk�exs>�y������y*��w��ԋ<7&�Z.k����J3)ޙ�\g;�@��	7�YR�v�u���1�1�{$�1���ne��9�?z�M����q �P��a��٭w�M�s6��:�R�-�a%BT��/k��V��J9��9��a��E#f���4ϓ!��������dU�ŒF��ilG����l�d�o#%�##"*�H6{�zJE�7�WN~{f���Y��v�T[QlJ��)������XЍQ�:)�=���
vFy�a`HMv� �/9��и�f����kTh� �8[H&kNF��7�R��"#��Z�Q��M]�R�C��%)o�7��6�J��yIr�e���M)S$����	��C\�,\͢q�8�f�5�0xH��CݒB�DЕ��M� �����E��(RT֠�=�5���IF�ZW���u��I�X�s��fI�9,*!C�&	���k[n��HP42����ؤ���	�a ��.e-vg���G�I���
gֵD/�\��$U�2�@2�XM�.X&����Q���'�"���<FI�o���|���}b�Y��k��Q�S���Ω;�J��ҙH�e#�:Y1�.-u{�7x�Ͽ̓�r�C�$`�:���x1"!�E� B��oUN�u�un���M�����=�眵|��F����(�O�و|�]7�Mnh����C��S^9�����6�Dn8���F/C����M��U�Y)�t33���@�InKR9���)���Ƌ��qtf#>��s� ��j
����-���S��e�O�t¼:nn+�69br�m��������������zk�}��ōO0i��s���0�n.C��0JM~�R
C�!�〗DT�.*�q�*1�u�)��D,��'`t�lT#�ʔ�[��|EH�	ʙ���m~�������ܢV�D�����S�]�2�EΎ��$N*�xF�e��l�2���c7"!������N�Y%AFgM�u����I�K�C�~5�ڱÄ2��3Hn��Z7I '6�[2��j���C��X}�����uu&1ڈ��pC�����mB)R��f�����~�s8�r�k60����Z�s�����34�rg}�:U�*���@�]c�"n(TD���:kd��0�D���Xa��sw6v	I��:"	�ѯ�)�j�1
�����c,2K�X,�s[_�]�q	�§�ђP1����Gb�u5]7�z�惿�+�V/��V%*�%f�J�5N9���j�{B쁄��!*E ֧��!�b�g��Ћ&(CЁ������s�(��g=x�"#:2�=#oYH�F�61:�8�K��}�ָ8p�>��@k�Z�L�?������hnB�P�P�׬+�1b篿�4�dn�C�>�DEs6\��OLJ�yr0��ϕ��3qiz������0n
��%�r�qr�t~�#|>�}�����]^xv?�*㩪�����L��H*.�~B)��Bb�	���;��e%�.CØ���!�!Q�����<�����O������	�ua3�0}��oR�*�(H��m������X�'N��u�}3�bR"Ā��۴:Z��K�hw+�5��5 �$"eJ2a�(AYP1{~��r�bXd����Sl�^��T"{�Ȭ���T
̔6�4L3�h�����l��f�j�!��:z�J)J������ڞz̡�^:���~���Ҭh��l��b�!��2%��y��%��i�VI�+��-:j�1�{�y�"��)�1�G�Y��(4l]w*��T���ᛜ��HZ!���$;ƣ��
�/(�~�e[1�	2��_c�%J$�rJ'��Ԣ�'D����%��TS��u_��!��� ��N�CB�ߓ��RYTЈ�PUD���*S!�!Z���� *��j ���XD��&j��K�c�H��d�L�<�1�c]��A^��-��o-�����t]!uõ~�}O}�z_J ��1�$F��AH)fE�����~�Zx�1 �gR�kI�u�<�q�N͑�I1�45Cף�&Y��T���^錒�	`���6d.D"7��i���.����fK�ĤP��nj%�&�p��^h�aYh�Z�y6wQ�6q�D��A��z:���F��S1�,�5��!��rJ�]Q�l�"Y�/�Hbێd$yT_���k���s��6���W�������$M{��j�]�|"5J���:���s�8?%:�|��0�yDFr��Vӳrg�Qˌ2259�1WsL�xҳP���Ƙ����6y��;�@�H��E)! �"!h�������Jal�x��Y�Ltf����QU�mkԐ#�iv�������Pe t!z���\��0�G���,0U"v5��I��}�����+�mC���go�R�����d�ߏ��nW#ObL�(�w;og��y����k�k���o�M��`l���Ҩ(������&E�!ԮÇ�4i��T���C�D?����֚b���l6��"HPJ#�*7Re�,�
y�$�T�i���prk�(��<v�rh�������diS�2R}��&w�
2����)d������
1�J�i*��&����$$� �Dw�f����uĠ����J�D�������@�2ԜB �
S"�q.�ɝ.s���-:D,*�\�c&/j�(�u5��CO
�ֵ�Ҹ�B�')O*����#�D�C�V�H�2�S
g�G�@`P�p*��P�e�ם�d�uF<���={f���܏39͢��1Wi!e�b�	�p��h�r��Sx�zh�kX���֘�3�
$��J��}l�&��g�랩�k
���I��э�=���=��2���STs����Q�{�HI{D�a�7NKa\��J����q(8��}�^���3`�p�6�h����6����v���X��'��6(]��e ����΢��|��ђ��7���@��t��&�2�\��ķ��w������!�hn��si��
CH��>�д�D!mrm����uE���dEP�z�����4Ld�B�p��U�^�h�1	�cfJ}��or3���LD^Dh #)��s�d{b*Fv�B��mn��ЛY�y�Ő
�f� ����P"^����4��
:�9��,�ѐ�s��6�E��t���vbr��*K�!)�$�c���\�dF-�R�R�����I��q��F�ژ��͝S�ƪ̸Oĉ<:"<�F��T���M�t)�w��bw�v���1� ��$�$���O9�w.7�!`#�T��ʦ�@[C�#ݢE\M�*�������=��&>@kjS�{hl��kL�U$�i4C���_,P��6�$B��K�29�<��$߳z��B��c�Qc��h���G2���u��C`A�.Bo�N���8�tͮӄh|t �nuB
�=1���c�w�I�+h	�xj%�*�7�k��E����;,�3d�#�`Bi�����[C喴CP�ڀ����j�!F�z���i�Z����ߧ�x	o-F:i�JVM	��E�J�aU�S���bn��W̜�iG��.L��1��[!W��(2ߧJ%�]N�뗷*������Ԛ�ύ#�Lه�U'Q[�w%M�c)�6?���m�M��9�Y"b5��
{���JJ���~��*B5��!D0��9GJ�{�h1�\�_|�}ϸ������K��ѫ�#4�]��J"S挕��AѸ;���9P�7 "t�==�4)	C*�D*�|�ǘ�̑[ހ�Ґ�ϐB��2a��06�Nl�Y�d����)Xg2�W��A�e8���;O\��i�BR �r=���ͽ�D'����Jg>KR�ds��=媌��y����#���J�@��<��L�֙�c�"��c4܀DGB��l�h��PSA
��Q��?�<L����ɐ��X�Mf�h�%/�uo��s6D������-���"�H��/oo�#K�����,��y�ں��!g�)�iJ�H��$ >�I�z�����7�P��Z(��������t�twM5�k�[w������xDd޼�B�neF�G�v�����o�A>,l�$�@�9d6{峠���4m�aCv��y�Xx�g���;b��RIRpő�GZ@�5̤:��D�9�z���h��m�)"_�c~Y`{`�GܔBz�e��P6���;nE��7>%�H�D��F��)�����H|ʢ�x��3������� Y��J�h�P�ќY|ķk-r(<��� ��-!xJ��ё_4�qCU�=�Uk%� F����HkZ�#���[�^q{3�/��.����Ԥ��isb����v���-�^���]�[(ۉ�)W"|�U�}�����̰4�-�i$�\���!G698h�0|�9��������o����
�b��hb�\^�xq�Sn��qqӈ�g���sڵ������0����'�q�k�����1S\�yze)=u�!���Ȁw#/\��K�*����$,)�j����fr�x�e����b�w�e��+_�ˑ���,ё�0���x�;˜��<�1��o��`j�]��ȩʹ;.�����������Ù�n�����T�i��j�z{sR�Ɗ��S�su��Z�{��<�?�&��Z��Ҝky�RC�g��Bk���rJ�����B�V�U���HA�-��e"��~9z�~k�r���;�KH�b"Iv�IH��U T����W�As]pN^*'��� X�3�pp�$!�c����i��=#��
N���n��A����o��d�6��qq$xSAg�qJ���nL�Z��@�1�;��R�E��F�
�����'l6[^�|AM��fC�2/�ݛ�>R�9�s+�)�\�tт�k�,goQ��aw���ܛ�������x�R��W�A�k���}޴�	�x�oo��M����w�
p�����%�4tH{�lܖw�H��/���Y!G�fƛun�Ҡ�֍>��Ѽ�kD��=��f�2/ٌ��3�܀.D��!�>�n���7H�q�a�3e�e#0�B��"�"4b7�a�m��������"Yf�)S�̜�"��&��`��֙�Ҙ6��7*�r�T�eF$��Orf9����Ss�r&�?�]Ct�Q�!nF
�Gz��M4�1ւK	�#�zT�W��w)�R2�m�o,_СB��$ZQ$��3��������\��������3�-2������?`���>f)%R^|��2ĉ�y��?��<�����:��[�af�|��F|���/^EG����_a��!U-�#c�Q|ʹV�!ס4D#18\�*��8�X]rl� ��y��R9�:��"��|�U_�(�qB^'���y}��"�_Qߝ��c����|�g��_�C�Q�]ù�k9���_�F��۩Z��'+�y�֓{h�ٹ֎@:g�ޜ*s�Öò���FJ3O]��r���՝uOϜ�*���um5D�=�̎<7���:���������	��.�brF�[7ǉy����A�k&�}�u�w�j��s=�n�3n'�i��I���Mu͜ǒ�ï%v̛C���.7�͎F#�D��1��g+gy���BKc)���:چS������ո�]�䤬�|=�(��3�BZPWy�C��C�s2�]�_�O'�$��Z(s�����!�BB&�|���iL̵�Ѧ��Ћ�����OD7 2P����J�P�z���VHe!��
87j��h�P$���/��1m�D�[ F#��T���    IDAT	��Dn�bMh���E������L��P������VR�OU�b(W(���TmK/+���H�̕���X��R�nwI	��%��&��C�.ʆ��%i�vxm��-���e�P�Ԗh� ���Z�aB�1�BKKG*-4c���Cpa1H��H�	�VQ*��@��q7%���L��}�U����[b�F쩞�+�.Ľ2��8��GG��7ҋ���-��)P�)��y$�Gj��WR�4������㎱���"D�\�]�)[>�)�eI0Y�t��[�ꩭ�'�PO�M�ZijUE'��� �>1��SϠ�պ9N��q�9���6�lzL���=Z�������A�)<�%����My���5݀�1ҧ�N�;�u���עG�-�Q�PjcɅ��	!,-����+.�#�%�4���5�U�Uzk8o�ٚ���9��8>��:��׻�}�ݹ?V��s���'x����V��¹�=��:��ʉ�֔���l4j�����ĸ��곟������};+�w��9!zo��#�O��o��> ���;O�c �礔�Rq]P�n];�NqZ	���:����y�����꽝�J�,����x�o�n�����E��ﻟ���kn�˶SU�}g�T"�e�FJNL�:P��/���#���yn�gi��-O��M���~�Ϟ�ɇ�Z;���>���Z���5J��e�Pm�hL�X���T����������}^�uq�\Q?����g����\�@+3��5�RQ-�h?Um/Z����L�y)�M�0È�ᘯlj� �F�Fi�3,�e��b��R
�9�!r؛d����G<��OUH����]�U���X�zp)��w�«��Ayu��E��z�W�َ�i$5G��h&p ^������ʡT��
��T�5�񔋷�~�>?z�){�:���ls�
at�1]sq���F���ea��7x�o������(Z�r�����}���{E�Q�b�LKPn������ȋt����)���{�ʳ�����p�A㊨�s煜�EM�YXJ�UJn��L�0:���L I�����
��c�&��	� :C�+�U�X	�o��O��G�Nܜ�Q板�� ��m��������F&����������܍�ײ�7��/�N6�絓��?"Ъ�P���*2z�*i)�l�;?Rj�u۸x�蒖�^='��pѥp{UwUݑ�sj�V�:�X����"���_c��z�{zIj8�3�o=�}A�j5��u��q�&z�s��wBc����^�4����e{91n��jқ�U��V�b�ά4+Dh�iՔ�L~ձ6 <q��b���4ܼx�&�cm�c��ݣB�����#�&w�a�=*�?�ͮ7��u�	_q�5���Kx}»�C7�(�����M�7���Ŀ�Ϲ��jtN����<U�ذ�-845<���<�����w�/~�?�*ף�4+���C䝿�ٽ�.���e`N��]QJB]�:׎�[4L�Lq`Qz��v�9>L�J����[��W����K˞��l2����o}��>Dj�%ze'���s"B�j�F߅>������HpxA���h��Z\@|o��:3ٙ`��^2�\�R������0m��|��9s)�.-�����[��R
�J������m��k��t[���W�%�W�B�n(M�U	"\u?��zN��
N�n���=>j�Lq�G.�/��Vn3�*'�~���}��I���q���o~�/��مK&��7|���:`���,�뛰q�q��7Ҿ�G��� 8�F�%��)�֘�t� �L���7y�?��y����Ң�:������p�X��w��+�5�0��G��r�� 4q�a0����$b�ɚx�U��R2�����hGL���9 ���~��Z
����E^Ϗ������j��Ί�5�iԳ^�E���79zf�T�:=_�;"���&�`�z�8��#���iv�Hn��m��U-�Ξ�*O�>bw5��7���{�2��):_S$�p�xG++��S���:^'��آ��������?�s�7Vhǈ��q�܃�wrV���=U��<�W�I�%��BΉw�{��������Y�S.�7P��}!U��T�lE<��~ֆ#�4������	Q� �;�G�=%��>)�!���z���GO����}�Ǒ���_�v�#��������}��I��v@s�J�&hT����O>���{�+���ɓo|��g����m��x�og���Ϙ��4t�
�%e�o^2uU( 7_��O���o�:���_%�n�-!񒋯�:�)r;�4�w ���	�0������/~��h�/q����\i��F.
^�ԛ������v���uF���Z3_�Rs&��͒H��s�f�.�E6W�}��|zq����r��Ƒ������[���0ni2�5<��׿_�����������,������ۏ?"�f}�=^��I�q���N��(8�|�W����xs���������?���Oٌ�O��?�w��=����?a�����B����=�����1�9CHz�"�p����S��~�g��IQ�(�.�|�?����������i1B�G��>o}���pK�����G�0Y޶�P����x�?����1n�8��Ѵ0��\3[<T�]�`�J,sk����Lo����"'��Y@�e�ۗmo����j3�k��}Dﾝh+
�@��tU��2������>� �ڀ�E^;\/�c:$;�9_��a"�b��^+(�[C-Q�~�)�.7�t@���?L;r9!+�Ѵ&�AZ�X�x$a�ms����A_�N�/��Ѯ�~挡oнX[�5��ЍT5(����|<�E�M�̫s]��4 θ��X�
�%F�)�<��f�#q��I�L����Z�b�xg]� ��'PR�a�i���_���rb�ݲO�DH��}k�H��cmP�������l��P��-�xh��{��&��]��O�5�v��'�}��e��8�r��ݔ�닽s��Q���	��y����:����bb��أ�!*��������-�s6n�&����T٤D�������x";.���Y� na��:�SBQ�af6&�)_o9��>��������pkI&ĒR�Cu�S~ә����(3��\w�^��C��VZP�-*���P]����1���CCD��=Sl��O��������a��o��ʾ��&K�'�����F��\T��b ���'�����ǟ�RX�5v^��5��	o��>n��Ⱥ�Z"��i8,�h������Hm�)N�Þ�����'\��_��o�� �N<_n�hQ_V��(Q��ָ#\nɢ�mA<qYx��������xk�m��_"9eR�ٹ����w@\FI��*�?�ea����f��J�����U6�3�J����*KɌ␢�������w+���p�v��o����/��k>��ȕ;j|��|�E��E��<��s��F�E�k�rV���~�_vS�U@E�;���=�
��ݘ��8������ȕR���еM�ٍ��˫--^|��z	p����F:)]�%{-��3�F��(V�z?�r�z���i�u1��qM8�U�;ό�EFZ֕�~�N���Dlpg5��g#"L����9�-we�@Ή���w�y��-^���9�^0�C�.��8!-�ی!�w�<�)ĥg^b8�����"�?���x}ҬZ��'�OTO��iP�ky�7E���׾�l�?��S,�����s>��u���5��1Kc)W���O����x��Ox���wx�k�3m�,@��=ڟG!���x���Il��!:�?WoF��5?���'W�3����]!�Q2Y3���,��q��X��������;/���J�$ejɔ%�<%�� Έ8�FX�a��E�L:�b�9�G��]#�ǉ��D��F�2pR��j��Ƹ��e�r�����0z؎�9]��G���O�oʿ��/�5�i��x�~a�3e/.w;�����>�	?������\����c.��f��?������������ʯ�|Çƅ	Ke��D�0N�\�B��ю9F��l�O���W�?�[�����!F�\癋�dyT*�ژ��SԓS%o_����Ł��=�'#�ӈ���ÿ�?���W�o�y�U"l`p�7J��ѳ�4�D�.hs8	��[J>0[|�hK�A�v��h*�=O�}����u>��}�;i�5�I��_*h=ٯ^vk��w�SQ�_�|?Ԕ�|��ߟ���C��E��At��u�ę=�oWZ������f����`eٲ��-�Nj:O�S�"JO?x�i]��;[_�����5���h)À��W7��y=KoT5R�6#n:'���(?~��]140��y��>�w���-���>p9�������c/C��h%�`ƢS'����V�)j'�̛�V�5B��8r��b5�*6��^={I:�<~t���1��W����ih�	s٩cP!:��XZe.��G�6��m�{OS[���>
�l��"�/.-�!�E�
�w��c��7����V�~����מM����U�fѹn��w/�*#��;1d��u>fΘ�j�pT6<�h0���O��ث��Z�Jw�:D}$"�{������u�a�w��rF����?�������6��:�w��Mp�)��W�q�e� �8����?��w����'vߝ���-���,�O8�k����Oqs�� �C�Ej�&�|��/^��~�?�S��5;/�[e��*������-���P�HnJr3��OY~�CBI��1z��}�������������4q��g<���PZ%�G��x�������w���e�x5|R^����?"�����Kc\f>��?�>�����?e���PB �"u#���*˼g(�����c^}������mD'�8�j�r�|�����m����&<�� ��:QO!�[b������߼ :����������s�����a٫��u>�昞σ��x�{��v��r���Dɉ&a���?���k���������	�y��+�hU��ߝ�V+������ǼD������������\\0��.sV޺�r��#���{&	��qB |������W~��x���L��w?����b��,V�� ��������\<�u��0j�H^0�1A�b�����4��E�+�f�	w���1��;ST�$���91���g�[�j�~��[���˓��6��]t� X��f'&����0�V��|iU8�5��(���a�h]����+���d��`:��N�DON�T*JN���%)�A�����Z�Gz�i|Ņ`���� ukYx3홮��P�Y�z�.2�ڎH�&��;����?�=�bd���n���{*��m%1��j�:Q��)�l
e1��������jI��z���ڼ*C���W�n7l7�J-������W�x�BʕڄF82E+�����&�i@���Z-�ܩM#]���*ռ���6���4uq�)��=��z$}>YW����'�yO臼�_�ٶ�����{��u��,�,°�Z%%�T���wb�J��Ȼ�}���1Ҷn�!.`B�]?V�x�KaօA�����_�����8d�y��%7M�8R��=cb�iK�,��U61 �X3q�si1�B 5�t��f������5�)sQq' ��S��(���9������ng�8q��v���gv.RnMhŗ��\s5�D��[�f��6�H�[s�������s�,��d�a���61��=��Q�j���1��)r�!2�	^�H�3p]�X*����
.7u��f`.��?��xZ�on��]�����Ы�������s��(�R��T9(���]�PepB�q@�,P+bPk����W��̣ݖy��4!>}�!0��㶨S������]PU�i��[�tA|�e�1��fp�Zx�٧l�:#Ū���s��3�՝9��o_�������U�Ug�j�.�������:��7�_�/߯�{mn�T �����~�~p��vF�[mO��;�:d�	�k+W�I��S`Z,��Mii,K1a�q@UXr6�,�0:6�@e��oQ�_g��FFM��L�	���ة�'�!@����e�xk������aI���g����WU���&܎�[r�a�q�����ɷ�A�Q�Q\��M��3�6��c�x��-^����3;�\�io����sF*�"�<H���4�7{Б���0��3iص�n[sW
RM>Z�l=���%0��'=��Rj:��é�u�p���qx�#?a,���]Ǟ;�g�����)Uz3�S����>����������{±;Y'#��y*�����m�|(�S����.Zz��)g)=2��W�c.��� <ǭz�ɤ�$
/�k��U϶A)�	{��L����˲�� �K��[kA��'Z �4mv�SE�.����".�V\̈́ D��4J�t�v>ࣃ Rf7\���=W�Hj��!��zIrJPpNy1?G/��fN�J����0�����@��ޖ�gCu�y8�]�h��oE�zOOp�Fz�1�4v�i�����)-�a�b�c��Ak?��nSX������	ڔ��F���]#93�A������g�l��H���V���yk��xo� XӡRL/�f�_��q�T	���p3^�U��a� b5�RjcS���9��J���_����f��glǑ�y���46�3L��U�c���%U�g��juV�r%���A	�	α�C� ޳Yc��NT�:�w>�Z�G����U�'�~O�9�:b|D����sJ��9�ֻ�q�z�ۂ��e�Ϊ�̓���vg�E�]�������}�riһ`�E>gs���ܹ�Cp��	%'��X5��`]�1:CT�RK� @N�Z*�
�������s��cٰ��=���ZMwv�>+=��}]�*�4����sZ���|�\ί�吾�ٓi���/hV㪱J��.L�棂
���͈� ��"�e�qL��0n�ˁ�"M��hT��\v��ֺr������K���e�b4A5�U���X�e�681��A{�n���F�������@����^���9Ϗ��w~��ϼy;}F��O8E���ؤ8r���Op��d��_e/�c�^�ڇ�j�	=�Ph��L4op�o�k
Zq�C�b��A �@��e�joQ���"�6�6f�v�z��di
��xP���ո �adlR��j��0������1�*�Ԁ�!�Hs!W��o�ugi.�&�ò�H\��O//�|򘋋�_|��g�y{@o
ZaOd)B��\�������@k	�-����D<T�/8�pq�0]�����8PT�(���Oog��	i���Q',%��#8�|)͛&�8��ni���E������qjg"\N�s�V�b��+sl��{4?�UJ&��s耶�G=���s�Ł�<дr��A�'8ӹo�����٘�gi����8���7b'y��RΙZ�aڒ��4E�0�X��1��09i����l�r�ŭ��� �j���9�����3��AY��F�}�N:�)nܩ���b0�O����<���8��Z��ޯ�k��d��q����\ɹ���@�f��^�Mb�Jo��x�j�S�TDgr��HK�ˎ8RZ���62āqp�m`��ymR8�b9����D����?�h\߂+�+��,���Ya�vl�Rm��Yg�v����6�9���x	(֜c㱽��"�8�:,��j���9�~k�pXP'l�-�9/�b�r�\g�����{H��eZ��_[E�������a��	�l�]Qs\�q!3�&���l����'��u�������z��oJ�2�}��|\}}���W�	�?�h�J��k>��5hQj5Czl%�J�6	�w���+�)�5���8m�
�*�C��`������8g�(��T7��"�W�bP.Gj��d�Z��t�-2'f���    IDAT3y6q@�#��S n��f?��B�F9�]]�|@T��JTK���@¢ޯ=��O^>�˟D]��-e� sZ�(ӆ�m&��f޳�'V�jR��&���xҾA�Vє!���%��X��U)s}����6S��؋3��0�@{.4e\U�`�JM�.\�RN�Ω��Hk#!'�Y�0��;Hw�E���cMK]�&\12(�fV*%%�'��<��z˱�v\� ���?x�(��"��2�%(5e\�h1���)�2�L�.�b�#Z�;T�;\���v��w�7m=X����[�����o��i�*�찵�6�G<-:v��K,�S�<��nk��ȞR�pJ&��q�P�d֏|���y���ˡ�ڀ�;u�)o�G����p�TH���HU)d\T�ad�N��U*�$���#�-�bך�FZ�qc�Er�l.6�&��7�
�zc7m�}bV���u�4����y\'�y͎S�3I�<�Z-8u�\Yk�b���>:�[����h7�[�"�Zŭ7�\��$���X��H�VZQ��1���`�V��.\ ���̤f�����a�`h���EI���B�!���Hˌ�B�ik�pJ&Yh���J1Q��������ܝ{�H)P}���{kj�o�ݽ�}�o��׶c��Ϝ��xY#�3퀳K���z��w�����k��BBt���`��<�f�;N	ZPi�V�-�Ur)��CD�G��s�}�s+4��8f\�N������s�i�r�J�vn��8ǒo{D`Q�2�~���aAZfF���H���$��QS��7g2�4��4�§?�!Yl��q��������?�q���~���L�3�ʜ��W\$�j��b��C���R�76[�^��.b;8��L��x��v��P���%%'�7��4��kj56�qHP��SJ~A<�������=L�g+օ_Gj.Х�+m��0 7@ȿD!�h���֖��-��G?��j��S:byr�-��т��8�r�H��3�w\��(�:PiH��2(.Ѣ'���J��i90��q�֮���E��������=�sڣ���=w��g�P�q~^+2�ϻ��-���(����|_��;)�A#՝��~Y@��vcus:���}�T1e���>FTzN>���＄R�W�l7#--����>YW�U����m�!�,kQ���ZYrb��w��R�䅚�UαJ�ZZw�]��Q��m^:�pvmb)_SM퍁��	�W��v���+
qN�f7@��g��9w��V�܌�c�<kj\��f��2]]�,ڼ���z^��������Nxh�����0db�a"�LM��U�I�ȃ*?�D�T��b��E-�r{3���v����z6�׬��w�u�ih�h��7}}��Np��d���A礗;З�>)~����s�sbײ2m��,�+le_���>�����+��w'
�!���e�؈	��m��`to�Xk��a�x�(���;�A���V�8��?G�Ԅ�y&h�hJ�>��0�TJ^:D�gd���^^�]#���!h@�����ь�?�F�2τM����F�]g~���=��h-
m���h��S�k�}�1��w����� �8�q2Ԥc����rN���q���G��K.�^��e!j#Dg"5��2�),�ď|thӖ༕��v$��8K���k����>�n�َ�Pg�Pc*[>z��\�Y�]#'��GU��l�=��X�K=N��~��0��=�#y9[��h�P���Gk!���j�~S-T�\1�$+��P��)�,� �5ѪJ�.��y���|h;j���������7U�#^u
H���u�����+���2@kK�:�x��O�s��:�IM�Zz��:��6(9�vߏ��Y�.=�݈Wؗ�;:P��׿#��*]�&k%�d ����M��񀋅���[��o������$�kn�ڬi��c�~�����C|��_�0=}������\i���N�%[+�O�Q�j���#��?�g�=��{_{������4�WiX�������u�jzT-�8�R3/�ox��i�>�M2�J��PGZ�Y�W"�ŎasA�������yb�-����w.ނa�fk��B]GQL�Mз�v/��@=w^����zop��v}�������C�{;�.x�5{�y����*Kz�@g��M��Vt@|�(�!���{AKD%��`_-��L?6rQnK%00� %�Zeh��|�<�ޛT3xV��]'_y��N�2&e�,,bęV+1�x7�RcVB�h���4��!ѡn`����$Q�ȸaPG)�P�8{�iDŴ�W���X�<syq��rxyMI�|���~�>zƷ�������	� �Ţ���P���Sa���V��ŅRl<��:�(2��sW����4��{�|�^��Uٵ�d�͞z�Y�b)�q(.8|sԔ�aKN�J#��8�[F�\W^�⬼`�B��*%-V��Fi�z)T��#c�||[�yyŲ�Bo�-����M�k#�r���%�K9�\���٫1����J���E �#�^)ޱێ��zs�v���і���~�m������z�����Νx7g�6Sz<��^0�w�Ȝ{�s����w�-��z<��J�ﾱڜc�y�.�T�� �.Xt�NΩX���q.���*��8F?ݡ�qxuC��!95�lL��nlڬ�M�/�VR��6��͋����0]�_|B���ޛ���6�t�Q_��B����Fz-�u��?�zU��7��y��'�~�7yY�j#/�.yY�W��6�d,'xwH:B��F�*����E�ӄje?�Q#�4�����u"`b^�V��(��0��r����Q���%�fK)��$�����z�KRŵf��5'j)8?��r���[oQUX��$��s͢U�Hp��E���Ur���4���@km��ޡ֠GE����9���s�HWW�
��ǽz�F\R�n�P�v�L/?A���=*�zB���x��9oz�8���=<��-�r�t�)u���jF��G��pp��/���E.����ʊ�X�#��Ѹ�F�u��I�z�zXZ5-�q2o�7{Quh�'��O]s�N:��aT}�T�kJp6~Jm��GA�^��{o[cG�����9mW*����Y�4T��1����霂+�$F/H5��&	_�3�,�T�����v�8	Q�y��l]�j�FFmf }0'Y\c�<~���x�Q���%�j�ʛ�8�:+}o�7��XR�g�k(�}����@��u]�>�4|���|H��)+�,�u��=��7bU��ֆ�@mJj�����q�&j��Gv��ԺPj��%o�n%��1�Q\��f]5;�fr̓B��:�B���X4'd��6�m\j�̅ZԪ��V��3���V��Yz�'g��k��f
d����N|��D�Jw̗k�V-'���kK�~1��u1d���`����~5R�u05�`����s\Q�ڃŪz$��J?7�B2ʺJU�if�,U�Kq�J�72���:��;��Q�$��{HD�lL�R�̭$kgެN~����XpZ�*s�0�ĳdX�FN�Gk��b���-���-������}�;c|Uh��w9+�zZu��h"V�OE��c��V�lc�9�.���^�������k����{��K��k�?�W�?�n��=cY.z�S7��NQ�����M{��F���׭r�����ݑ❩�Փ>�8kLc�F���^ZY�䃋�10ω�^����l64g��;謹`�g�!�V3�v]ET+/�x�n��bsII�r�hCo�lQmNq��a����a%��^�A���m��:�	sꝰ��t���|��2���&݀��9�2�z�9�'︡mL���=1՛f�H�qk�%��ȱ�c���q�w9G�1!"0"$�t7�����;'#+�r�iV���5b�wMq'�C� A��w��Ĥu��7��Y�أ��S�j�~Z�t��=,5��j�-�n��Js�1R5� V֔F�LS�������'B` W��L�x�n�����'�Θ�k%�)j3&z3z��VL�C:򲖺�g���,���H���Nc�����.�TT��+9�`ZQ�K���*9�B�}l*J]y0!�HK���;�sj�j�^k�u�'�%:Rͪ�#�(5���硘��e��;�\�_�)~p�spǱo��5��9��U�lf{�C�Վ�{H��t�ֻ$�AFkJ����br�ꏟYsˆ�YY�ݿ���~ޭ{����_`w��=0�YNc{��|����)���`�Ɏ_�e�gh`kJ��;Q�mp�*h�߮C얶�t�6�zq��9�����1m" ��g�{�N�qv���v�e�F!��q�۱"y��iDs�c����}UTtm�R*�+-J��u!_����1��b6�������������O?���o�����<�֬N�9�T��u%(p&M{m7������8�m$l7��k1o�K/&E{��0:Gk��
��3�er�y꒸�3�43��q�@�4餌��3G%�LI���������C���Wpո��t�����͖$I�,�ò�����K-�C� x���?��'D��Y�����r	_�Tea<0���gv[QT�{������r����f�r���D�QD�a0"v�<�7XN�4uF��G��s�]�,�a��3��؄�����0��ݔ�k�.�0!s��d�6�7�E�aF;�os�mJ��!��x��x����Y*�[A8�:w����A�6�)h3�;�9`�:	F��(����hmN���!�qs��e�f��D�hChD�-6tE���g���`G��\��l�U��2nD�tj���j���ϧ���LZ.<�7�Q+��P����O���3JJFT��ٴ6Le�����Cbk9H�0�]7[<�Y*�V�.�3��5�P�������tla�rX:����1�^�}'���q(;�Ӑ��о�sv���ș�c+9�ّ�w>K
����tO��^�ۼ]d�1�1L��0��Â��bF��_{2>��On��c�Rb6K���||9�J��P-F 9�_�,��MG>�e��TH�C�E��6$��}0J��H��YmJqTN���yA9��>?`�#�D|�g��;�ZWX�v�X�I1bb�Jc	�l�S�
�b�u��f���Tn�jľnI��(��MEv�.�xX��{��s?sh��S����^����Ϟ��`ju�VU�Py686��r�ũpN'T:�զȝÅx9����[�f�Sz78�/�&�ղ�1��l��Ư?�J{��p���P��%�	��C ^"�wR4(���l����,�[��t����I�Rv��Á��2ڐ��lm�0=Z�t�#�ﵫ�C�`�9����#"�4X���x�����2O��%3+�kY�<�P�)���Yt
NZi� L��}�Le��Y�p"c���߬���i�j��{T�k�cb��"��jrF��_��b7�A�
 4C_��6RA�VgAV`<?���i� ؤ�ٔ����a���6��Z��5�ua�y?F�ʆRt!uA�r�"���&h�ZPQ�����<���]��P���OI@�?��Ð�!b,�ʡ�{G5�-M&��6Ku�T	�S�I��G���ű|XU��Y����րgl�	7arg�sl�!.gk�G��~�NA�q�FW����I�������X����Nn��!�r8Q ޟS{�5X����ƙ�e�|� �m�:���;ym�8�������yV�!�r�9L��k �2h��ż����)6| ����ʆz�=�s�t�ْ@Z���1G�j��h�!��*�*��Ļ��#��}]ꊄF��]��c�B�V��Vj�x&���s�!/���Q���l
lu�|Tk�%�#�V��#!�m���y	<?=Үo3���G0��xE9��m1ӵ�$�8���eA%�$�U�f�a��xM�(L��ӪKbm7�m��L�'�U��T�0���Zk'�Ľ4�
�T#�kᵿ!����m�vc+�pT3 )%P^#!X}��n�J�V�����r��/������1�����Go�6���V�3���B���o�Qê��C����!F�!�5n����\�&$�[��jd���Ȃ;z(���y��o�@�l�`�|��X�a�t�X#23*m{]2�.%������0���b������2 ��CH,9[�Y���2���$>>y�{���F�Y<�R�	h��`�m��MYͥ|{G��x��d���#�<���r���'B�kߪ9��Ս[]Ms"X~SS����һ�I�͠X�!�N�@��J���H��G�������[����9vOI�s�_pg���"##���c�$�>P8�3Q�\i��@s��9�lpk3�f�2�����d�iI�#��FRFZyAe��wvR���Xo��O� ���°rV��,������"l����s�e��3��{ޯ��(S(,ؒ��,8~����D���Y����Ltڮ���9sQ��}"b�i�f#�kb0/�k!F��6g&��!
!e�5�uk+-M�7�SB{#�Amo��I�}�p]�NeSj)h��xך=i<=�8�DVE����9m��3��)h�Z5boy��]N�P�(�%�P��bS��\�߇5�A>�T2�J RK�u{'�L�����<���g�t���+���9�0���0�s��˼�b�\���������g��3��Wֺ%�b��&�����(�j�F�H�Z�K�n��^�<~��~yk;[y�ݴ��Zc
���1U>핪cSF��Vjm<>>��Bo�u�lxdM��'�N�.#imdGf���GԦ�FVs�k#���>�HH�����~#�;�S�&�q��� &$��饅���%}��f�]�V7� �h<�m��:��tmwL�m����`&�:!]i��Õ��%���1Su�X�1R5g��u
&�;W&s:�T}�T�g?��G����a@����C��[5ti�-2��CF&�N��Mے��m!�k�Y��;	r&�Ŝ�w������+�?���_���C�c�ڛ%c��f��j������<�8?d$)�(*�X;�{�@ӌE�m��0z���պ���Gg�q�xO�(�L����J��Q��ڇ��{�Q܄MR̐��v��y����:������]`�~���Ӻ�{��M��3v?��}Ԕ� pu���@����!�N��0Y�Q��|8��r�mT�3�UwP�!8�'��x��)3`i�{堾vD"�����9�E�H��¡R뎌�fm��gQ5��![ 1����3)/�/���l�7�k�68��F��ɤM��Z�8��Vr��(��R6���bB0�����D�{Ta+����� ���Y)�"<=^XN�V�`��Z-p�ބ��^�{o�38P!$n�Fi�ǧϟ��]���<`�t��'K��g���gIHİXoj������������G�T֯o���D�c���B�&#�gs���ڭQ��x&�X6�5���߾�ť����G�j�f8A��bX8��`�u���-�(E�����M�l�p�V��ƨ{M#26h803c���9�U������R�A�}�6G�96\�m���ё�F�N�IL���
ֲ�R&�lY?5cd������s�i�g��8|7/���,�gG���d)��[?)h�A��t���0
Q��u�V�ɨ{�5����Pw6�Tzx���0�ʘ��{wiQwnU;9�C�:X��ޯ{m��.�L�'��˯|~~���o��o�o��������`�w-�u��.���R$=���;KH�Ţ{6���dpd�56t��ϟIKFc0� �io��� �N~�Z���؇��0�!��W9��a�,����Hk$�,�;�iPH)��Q�	�@;� ���q�6��r:�{���N�vuv����n6�.I ]N�� �)�H��h����e�r�;E��y��t���=ɚ���m�F�s�N�����6����k��T���X"a$�Rl�n��@�<��ўqe%^�ۥАIO�.�<>���|���'����%���j��RM���&ք����e� �ZnV�	�%�{��a��8ؐ��J�
�b��    IDAT$�Y"�,��!r~t��mu1,�[�n	!�I��[�ݻ�$k��-q�*�N'��|����(�+�13S�Ds̋U��9�5VH��C�P�
����	io�7�ߕ�ϟ�<<�����u.��U�"	�^Meo���T� \�k�xy�j��w�9]N����q��Y�N�7��m&	l��(��4�S`Y���X����\Ng�uֺAJ����DR
�`�؜9�zb+7T!�̦j����xk[ K����3y[�`�CF�kxK�#_��l-��X�f�lP!m#=26w.��k���^&�AV�uj�o-*$C2,Sj��`1+yl�L������|8���(M������'�vf2�`�1ͮ�ḅ{7P�:�1���%;�i��H�YT�p��w���h�&��s���u��@�p�/���D[�+uNt�5��HZ��`��A���t��;_^.���?|���﨏gn������m+��+�V��,%���/OloBt���ݨ��$�L��Rh�wٚ�C���&��&i	�4�
d�!)JU�]u�U��10�F�9'|m��HM��JL�H�<�j��~ə�[�3�Q�d�4�.�W��B��L{ ��g�${0�?ޚ%b���{�J4$`+j#�P��%z�L�]��R_2"V�Ӯ�_㰣��@��=���;�ټ��&Ԁ����f)K�3,��3끎��%�s�ڏ�����v 2����1#����1E9�����V0�z
6��K�]��pyB���e}54gb?g�VC�:�u�6�͏6A����ҭR�:��=��\i}�9&2;0r�<Ӫr����b�pX�]@	���T3$I���2�Vu^R���
)�ty&�2o�_Y�_�a���K=�0��Qnt��@xRj�V9W.�;Y���������w<�����Ͽp����<c�	hS%
'J�,��(j�����ˊ�;��.���򕗷W.�D\2�m���@��
�P{�U�jxDͼ��~�<}~��r{�Z�&������X�g۬�r	FH���46|�$�j-b���#H!j��Y&�j��Ƣb���B���N���r�!�en�	�� �Ӵ��e�p�u��R�7-�V3r�6�귮��I�`G?�WwK�����8a)r̬ňJ!����s����$���?d"�B1ط�|�q��%˖T���>�Lǃ'�5�ҝ�m/6-�3�`s�1���N���m��u�(q��c�ؖ�8	RU	z�`��Wv?B��Io�*��G�s����׿L�\{g��V;�(��fk+<=��ӟ�˧�Vn�z�CR��b��v-�Zhו��2�l�nׯ��g�$&:��- %�I�[$�i��"��F� ���� `풃+�X���/���Κ?d�f�0�1T�D�+J��m�f�2�ZmνT��9��h�
!�6���}Q�z�(�hF�=����+m<����]!iY���)�u#��|D|�Z�d���$Z��2�N�MC��E%�H����:�Hi�#�$�}2fp{P)�:�g?��8:c���?�J�A�T}p���^Wyk����=)-�A�@�yy���5�Nc9�(
��9}V/������/?�7����e}{���Fh��9�8�.n׺�i�����$7bwm{C	R����nW�JΙ�t�z�x��+�2�l?���?��?���o����k-�,�P<�:�jc�<�z��}��@����n������K�կ|���I!�MuT������UE����M�ZY�:s������*i�MWգ���yV�^ot�ʷ�~AKA׫9b��U�#�32�P���j�e}���x~�p9?�B��ol^O=�4�P[&~�K;�#�4��0x1���ە�ϟyz<���B�m�:`2[���T�����@��u|��00i���:ؐaŻ�4
O���)e���|:���ҕ^�y@f[�ȆB���(E{��ӲCkGx��ꆮ���!��a��e�ӿt:�CՆ��f0���b$�LΙ[�~w���ۡ��N?%���u������$�}��l}
��֦�*����>Iy@�@��ݏ���r�1�9���y���2|�?�2�c|����!h�#��,�)Gj���:��������o��+�Z֊�kkH��QLV��]���iaK^�ˬj�\�wB�.jYM	Ѓ��=�7��1�h<��J�1���{��?@A(u�HY��u��9����{���!��\JJ��,�C�9��l}��jG���M,@�vӎ�u�� \�z-�%��Q���t"�ض��%��N����I�m	��l^kC�<��Bi;5׻1ޣڜ�.�×m�7�T��ujܗ�#'ALJ�C�nV������z��;����9_j͈�x� IvP��W�G�d6�����1r[�����\�ty&���yp.�	iS��Ѫ���H9��[%�q�8�h{-@�eYP	\o�+1ejSd����y���;Nb|������:KcoOrg0n����u�b��'���@�t-�fNKF4�B),�]S��q�:V�#Z��aU����B�!ok�!Lݮ+���t:�������+/?��C��by�q��qw��&흹r��x�+��J�����'^y����Emԡ�'�.�,z��'.|�Չk���)+'�Eٶw�m���n��Ƕ����{���QBV�6�d�pc�����8���D�"��d�񕸊���P�0rb�� q���&!L>°���޷�t�jd��|�0F���z�!�?3��2��<���̐���>6��׮d0!̭(U+�6+u�3�k^�/���wcī��Af+�(�$w��c��Ww8wC��襶a)ѻT�~�L��u�AΔ�TTrlB��Ht��G?KL�^ho_�b���ĈS�F'��rC$��ڄ[��&��BdM҅#�K�9=����9�6�Qa���@8eB�4Bs�'�}ks��AN�#'��urwF3��A����~m#!�'�뷯7%#�T3A����/�NB`{�3j�Os�2$+i>İ���#�G����~}�����	��f�KϾ�G��?"�wO~��=�#�����C����#S��dw��CJd����n�*�b�ǘ�v|&��8"b����[��Ֆ-��N�u��n@'�@:_L����ƞH1�{��B��3E�����I����*�c2ތڐ���Z"��eI,y�ڽ]?�%PC� B<Qk��v�	q���mE����_�������J�@P�8����:?���V�J�T��{$ʒ���Ј��7��F�}�Lm2"M�����9q�q�0A �ԡQ[�/�ÛV#����?��G���[����Znܮ+�6�Zͣ����$b���쯷����S>�{���"�����bo-���6c����L�ǚW�ڵv�ؤX�J�6��_ޑ�<>-�4n�m��¾aǵ+���g�J?԰�����{��2�1��_�V4�嶡���N�9���=��n�ʣ�ѱO֟�ޫm_���N�u�����ٟ�m�h�o2�0�`�b:H��EH)z���h�h0�r�����b����><��48���ӘK�%���?1줿���}��C��Mb���!HQt��}E��$k��K��Ih>�����A4Cjm���|��Z�Uʆ�319z}؟ɾ�bd-�m-t�HNTU{FR�������O�vEk�5����^^DWNQ	�����pS�m����p!xy'�D֣F�DW��4��
����Q=�>"lл����Ő�Z������2Z��J1F�)s?��Y�F����~��,��Hc6���'�yю���Q;yQrzv��Ze&a�8�l��� ?�r:r>v��\�[CEI�I�Y�$H!�5%w{);��sH� f��	DB���9������`c�h?
�}�!]�2�Y��"�$'��4��|�dR�p�Po$:� ňF��Qӑ���dZ*�7Z��1��uR�=8K��f��*�������w�|��rb{}�����ѣ)��n~a�r�l�l�Q�fmv]i�WL{Ɂ�ǅm�L�w�Z�i$�W�CV�8�L�:u-��M��KB��H:t)�*4j�:���S��o��/���|���ߨ[%��Z�94a,���C$�`�f���$Z+\�WZU�ϙ��GzXY��M�\_~��.��;j���U��DA���U�@N�N~��{�a<��қ����-���(�ea�A� `�8Vֳ^k�K�ݩ�f-!ð��򏤔�X�r�dfV��%�����Q	����&$Hw�+x���	a�;f�m��wZu��B�_;
>�l�ɸ.q�7#�Egm�|n�_�}���D�!�~��}�����������[8֣�����bm��v�P�3�H
�NQ��0`�����QkUT�!��l��o�f�`��O�
��7nk#��UZ3����O<��|���+�ۛ�y�S�d�:d�]�x[�Ѵ]o���4'���8�c��G����S��?k�s�8?�� �������+0v�Wk��A����e1}��5�d:{���:�]��?�H��6�N�n�f0>��u`W?�`���K�� �:��=P� u���Yd�>GCzԵ �;����A��!�8�/���{t߽N(����fɦ��]Iq'�R���7��?/��{��&�-��1�h���J�m�vEz1�J����l$��yp1�AE�O�쉃�V"1g������H��VMlkY��'.��������#)/;qu�w�
mu�֩�ћ4��J���x��f�wQ'�=�ޫ���5����'��]����QSM�����nd��t���_~���O����}}���?󰜦$�� *iD)��K+�E+)�ڸ^oT)|���|1g)��Y�E�^Gq��7��?J3Gc�>�9�2[]�����8e���)%9 BT�;����5k�È��'t9(C��y���a��Ǆ}j���۫xvl�ў6����`������uO�-�5�q_U�*��m6����g�c��x� �F�c[�)�)0t�9
"�όu�����j��"�)@��X�����b�7��yL�Sݯ�~�������7��3��qY��uܯ�����]�~x9���5b[�c�[��ڽRZ�Uw"�3�`��ef���7n׊��,��7�=�#��+�me���a��ݠ���j�پ5x_)Z���Dw���$�N3pb�w\�N�_�����ZU���͞������d��%��;�`�@�	�	���oc�Y�%:Y�Z/G���`�RF����6��[�J5q0���S�	�^Z�l��r@�ܴ�}r�C˲LG3����ahb����c9
�xA��/D���2h(���o����	 ^B�62����1}���9yڑ�n��ZV�"q$5`2ϊ+�Q�T2lU�;�Ǆt���v��g,�@���rZ8ga}1�L荭T�c1z��y��z'������]ń��S�$�Q�-�s�&p����1DZU�V�CJ�*��?P��J�Z�?�99t����K��"�/��3O�?�^i1�_oj�g�]Q�֟���x{y�tY���"��X^?��=G� �nm�5XF�=�^5Rk���P�V;J���i��8�hl�!�c��Z�v��GAw�s<(��7�I$FXٶ�M�9�%��l��U�.zW�7��9�ׅǿ�u������-��;:ϱ��2HJ�|<��i�f��p��w��x�w��k�J� u4�>��]��}���P-�1�:����xDo�׼�h�����(�=G/�1�<~-������%�������>݈gA��]��y�]�TV���˕�늰b����9/�.�����L�X�vۨ[!���|F{3d^��ͅN�
�y
9�il�}O�L�u������w�+ԚM����m��UXNy�B!�Cz���]��m��7�HG��cV4�1C�]���K@��NPk4���@$	�X#sRz���ή�[�>���s�>���%2��D���<c�W�h�e�"�-��F�5ǿ{7�E4v��|BD&1�R� Ot>Q
5Y犨��Q��G�j�w(���zc*<��O�%H���R=�:���fB����e�S�JJZ"!��XWC��u-�R�)�%P��΅����D��D�nY����~�v�,��I0ښ���J���]+�����4$$䠼�����z�"��~���[W����������'���o���<�B�$����`���,KF�ZP�I]y���V�<|~Dc"D3Z
��F���,\��I"J�+!$.�g�Rx���`N��#0�@Uw��y�d8!�y�3�`~��У�hJ�������Q��V��S��#�#�3�>�Y��d�z�^�!��a�����:�ޒZ�h8�����d�Zf@#>QK���#�=�ufo�M�/�L|�=�p/A�h�[�u��p��!��	199��m�D4<�W��C�~_k��J��r�x_����弣}�׏W��}�_��L�����S_��6��3"9�]Kq��3�X�7������ڔ����oN<<,���w���+��|�Y�1����SS���P�2)���ϡ�w�X��TADfr�}> ,1�LD*E}η�ѽ<d�y7���q �F�#0�=?��u�8����j�}� Dw4Sݔ��$��z%�L�f�SJe]iZ��i��Y�e��-Xѧ�uߓǵ�`�(����zi����˾�m��1�c�
�y�ﷻC��ج��6�A�~O9y�����8�7Ė&�ب��l��$I�s��uݸ�������������b(��!�q��x��u"�3`�&��Z��F��O��Lk���NZ`y8�{!4!&+7�W#=^҅Z:ۺB����jU�$��\�3/�e��2����Y�Lal�	��`��ڭ�q��n�>�g�=�N��G�1ҥ�����]��ң���[����Z)B����?�H������?Q�o\b�l~|��xZ�(���\΁��ޡ�B)J�
E�|y�v������c��?�ȵ���ӟ��V��
����6BL,Kr�/駽�uc	���k%����'$(��;Z*KJ�+�OuD��s��>X����pt���Q�U�^��K����C�k<��"���Y�ץG?�^K�9�:�xVb�O3��s<�Of5G��^�m ��B�H��Ԁ^��7m�nP���f2�D��N8��K���|R��% ��H�atyxPq2��JoJۜ�%m��)����=��V���0a���|O�n��x{��4�bD���N�]}mώB$�u:��7����;�y�d�Rw�0����6V  c=�h�L��b�ڐ���r@$�5КP���v��L���BJ�?~��C����-c�sMV���{)�����-s�AL��k�q���Yׁ	�`܊ �f�+���ZY�d)mz�u%	H� �7E;��:[���rds~K���h�h�l��[��A=�n�v�F�kx�U1XKcS�H�{;��
F`s2�`j{���=���w�Yvfw�Ӏ��	�!A���ҽc��,I%��i���>_}�cx�������Zg���}?!�b�	�i��iN~k�ln�**c�dDz�D�-(�ۍ��ڸtK��-�q�]������ၲ�}x�&��wD�9R1�f)�ꉘ;�����7>}~���L�7�f�|�a�a5�&������*�n��j��9/�/���?}��p�l�7��J
�bø���V�t,h�r���q[o�\�
��d����Ø�فt���ul
�`���9:�������3_�u�U���zv�V��w��#�=33��~��S�v��+��~���������Dw-a�g����D����%��x���[m<}zd�<������=UBP$��Q��e���k�T�=�-c�3u�~2([��	[��>�9�N\[����m=}߸$�0���d�"�Q}����\?"-�Hv�l�&�ʄ���ߐ�5�I�� �H�;��2�h���o6��S72V��,Q����輕�$$sr��0.n蝗�A����    IDAT��I"$��ǭGK#8��J�;�4j3�S#��Z��c϶��n�gf�%W�Sۛ�Q��X�/s�a�3������3���T;co��l�鬊�h����i~���V�A��(l��k�r�X�p�7�3.u%�dħާQ�4���e�C���8M���nZ-���&q'�Z7��u�3��8��!����0���`p�RZA�^F��'2���=#�4|�3oC���q���a'�^�ξ���v�^�z�;�&���`�a�Z�ҍ�-n���A�e'��%���f�(����`鼽�k:��]I��s̀�k�>V�W�l��RJ&��>?}�l�>�/�bk>Q�fȡ�E��sF�u�T�&�M�.�͛�Bp�/�Z��,S�\�|��1����.:���l��~�g;Z�)�ZXNg�e!'��
]I�H7�+I��p��s�)�,��f0!��6����`���Uc�t�G�	�Q�U��s��Y�]鵑�|�-����__x�<	����[��^��Ն�e�����;�$��|�����Q�-�qm3�2\�`�t�����wd���z�Мy|~��N�+��A"��?�3��]������gYz�� ����*g2I"/t�3eI"9�X�HA�{;D�|x_���3��<��ؐ�9�w���0�A�vG�4��ݟ���Mb����g�DF����Yk���i��.�@�τ�8~���+1'��4��g��bZ��L�`�Xrk��]]�{G$�/�n� �(2�َ�c�l���|]\ip	�5���������;̯�\�5b��Cj5Qmʲ,ܶ��Ҫi3�i����e��%��U��*A�_�_׈�FU�s��=���S�^��LUd�`�3�1४����$�V�\u�������n�h�����F�{3"���A!�*����9A�퇝ѵ���3����^�ׅS^�V�<8? �H]]�  @߿a<��^�*�L���:�r�GX~�hZ���}T��¾�K�k$�Y���׬���S�Mq>@�Η:Q��������^��2a���������^��k�q^N�[x����a��啯������LB<@��D�q������V����FP{	  �ħ�.���e��W���I.�����Ȯ�C���%��޹����Lk�׫�MF��^���>��l���/�Zk2Ѷ������o[�g�Z��<��YO��F:������(R_}�������E���F�B�HjX~���6\������UDx8?�^7~��|���6"|�O�D��T7�Zw�������t:APޮ］���Ͽr>�����d�`���-��V��p�Y�f���rZ��*���p"??qZ�z���/�/۾�F	a|^��Imc��Gtg������:��M�Z#��ǽ;���/���A�k��6�=:��[��5�����ĸ�����됗9io���+b7�{@ћ��6y���k8����b:����3ه���C����!֨VO<>�=(�A2���GC%b`K����R
1V����6�5�9�H��ƼJ'����v��&Fܳ1A�@U�Ho���BV6�p�������w��<b�l����INRӭ�e���?]��x˲��j���9*7���m ��l$�pª���X��`������h� %��
�p�vV/ըrzx�[�c���n?ND����|2����}��y���N�ϢO�I��0�p�Κ�0�f�0���U���T����`�n��;_1g�@o�{k׵��kCc2��d��O����f���A"v�B��y����b�$�T���D/��	Z|t�F49WB��aa�����u]A�eݭ{�݃"\�v��ɘ�>�z��6HRi���j�4�RU�KR�Կ�H��J��h3v������=Ϩ��㐢4��H2���F�]tv��S��ps!�#G����_~���g~����������������#�wX-D!�E�CY�Ғ�n�_��\�dI�r�Q����鬆�!�����;,Փ�m7�V���(��(*d}��Z�+��vPN�h��^>@:D`gzkP�j,�rY(�����_џ����¡�[}]j��gVÝ!<:�;"B�23$a;��߷�Hi���A��Z��ѻ�RӾ>���	Q�wNN���څ�;2�ӴڨIsZF,��GpG��+��uOC�3
�����['<�.��ZvV=:`����s*�����;��C&��)Z�2�q��3�y��47P��8#(����S�k%J��a�i�����y�~�*F
�.��
�L\�H)��I�i��v�b����B������w��?G��!��;7GQRJ��8P$�j^��hm�ᔧ���X_�۔o���q����s6�|��g��8��7k��F����)-���r8��n��"���D[� �Uֻ�0�a�析��6A3��2��F,�~�Xy.��c ��(B�*KL� 6�v��xpU�k��aذqԿ��7>ܨR���K����<�U �m�Sz���3�6�v;���c�ja��})6L�SI�>0����l���eA���M|ʥ�k�Ɏ3�H��/�%�M͡�à��1[�ڍ����Ҫ�Q)$Z�.kl���Y���QK!���E�� ��B�C���ԑ��LAМ����Q��xGֿ�3j�'r�JrSʶ�ӏ���~����o7�bSԬ>b3����4��Z���@��^���tJ,�رe�h݈6ֺ00����na�ť4B�콭�A� -/6H���Z����d��9�Ȟ千�"�t^���k�\�;�/_�[�tna�����89Aj�Uv�������Y�/Af���,}�u�kǫ�6K�{�g>��N��z�����5���p5kw\OW%�Ӥl�Z��0�"wJ^{f=�F'*`�;�`d���3�%���#u5����q�J"�41i���i��8���=�m('K{��[��l�AN�4�;5쥶��Fk#7�s�b<G.�<�ǅ�ܱ�T��>�ӷzSn��ֆH��/?S��0	b)(�tD;װ�e����R
�2嬏�mH���v��Ht���P��5c4SGi)�Uϰ�fS�؝��q�?��~l3;��"�69L۶�sO��&?S��Ύ�֨�fA�����@Wb���\�eڞ)��{�?h�����sj�'�h���j�Nc�`�O��έ}k�q��}��P�}F��⼗�*9��e�L�uz+N��D5R$X�BZ��_o�pqG_�������N����\�� ��]�= j��9���E|ts���9/3��i��1�r�i�k���-˞-�K���I�Ր�$$i�!d=@�hC�<h��W�SL�٣�{��V������il���![�zP:��|o{bw�^���!U�S>�믯�T�� >?��VL���J�3��c!�\cX%�-�[��ן�r>/<<�Y�b�\[��<�#�$b���Z{UJ#������t"/��W�Ĝ����\���}�}�t��L5s��)M��V7+Ah�QK�Xi��}fXx��g*b��J��Qug�Ў2���~9 �Q�7�]6�$DuE0'Z���&B��X�Bpy�N\N��n̋G-�4	ʽ�aY&�H�FC�9�4�&J������Yl0".ż��G�02����T� B��=Tw4�`5�#
��I�\������s98�Ee�o�޾�lzyd��ܣ��KqA�`�(�x����GT;����,��}��κ6ҡ5�9+�J54oIg���t�:v�z��B�2,��f.��l�J"Y�hO�:5�[��1O�����ԞY�W��FJYm�e��;�@ݶn#X3�Y����zQ��[��<g+MY��ȠBo��ֆRg@�u`��0�g�:kԣ�t��K+����!�q�TJ��:;DDLR{��;ik|Oș�d�����n$�^����"u�h�B�ɘ���5=��y^V�����4u^�)���n7N1Y_	Uk\oW�yr}"6V���^lVAU%���4���f�坓ٱx2M�L�ցa�Ķ��Q�ּ��B�󬝜")ڌ��6p�	\
؉��9'����R�)�FL�6@,�A:6�3��D����;����F�jD7=��.ku>�mL���&d#1�Z��ۭ�׿��?��|��?�O��O\�!���% ��@����.�%Qk�VV���E���J!��%&na3pq�z���y?������9/k{�B̰��(��}�����жAh2���G�@�t]	�衡��SK·0��L���Уպ��d����#z��^�;�U��d�0��!R�Ü~^>�jR��$Z�S�����աe���3�p�D(������j(e�Q��b�1�LQ�]M�p�66S=��y����u�C��w�߫��Z=���~#�0z��.���g�2?{8i�^�����OZ�ȪF���=^f�=qØƔ�v1e�R���ӗ'BR���ϰ^I!�$�4D��@�UM�3ҺO��H�M7�����<�P�ol/?C/���I��5�~eY��i�氆������׶��e5�Pk�t6������|��qi�;�Ү%�ĭW#�a��:	2��w'G�����>���Ge����9	37�큅H���a��wz980��!�e���U�-˂4�>�� �mx˲x7F��in�F��n�{H��Ό>i%��6r�7J�{��׽�6�Y�1��O�e�^ۼf���6r�lj6o����v���˅�9���t���#����%�l��8m�%�}�1@JP7z�R׫�L�	�]Ap:��Z�Փ���m#ˠwg��ɫ'5~�G���j�v{'�|X[3E�~N���ڶ�x�<��2ݕ�ɞҴ�j3����H�g>.�����]_����oj<��72MZ?x��,��x���2��x��o>�W~�翐_7�I��N["[P���x�βN3��PG�&����Q�jᶮ<������i�喻~�{�CD<
����5�mv���OG�;��k���9ϻϐ���1�5�߼?B�{����3Q��~��qݎ���>�&+����ƻ��l��q����>�����?=���T�ϻ�\�S>L���k<���=4���a�!��{�G�q�����b�!����ܴ�c"���J/I��pjgm7�ϴy}Y}ȐA�M�Z�ߞ����?��t��忠?��)�������˲p�^)�F&�Y�E)e������̈���gdJL� [��W�ca:�a���3ݏ�������<y��d`��}ODf?����g�[{��(�$C�B?��k0+��؃���ẏ{k�ϭ��ڏ\��a?�����"=���L~o-��ͣ��?�O;�x|�]{��?7��du��B��s�RʨD��>%1��"b×���7��I�#9z�NFDfuUW�����d�+���.��J�Ƥ���~eefIw@? �;�=˶�̌�8����"'�0��J�aC�U��:s���)��� C���:�C��j�prb���o��������?�#菲'(�Ɯ;lh۠Ù�Z�������ݰRN���l�۲`΄RuY1���~Ǒ��!�Q�.�q>]p:���� ju�юQ� d(&�����pfz#OP6�.��~�5��ѭc8��ѡ��y�܌c��Z��3������g�����Ľ��Q�B[����$Pk"�{B�Vp���?ˤ~4f��֡��x�ج���5r�V��� +����I���8�Z�c�}����Vm��p��lM�8����P�XS�m]�{��iB�Q��� �mi 3�|����O�p�rF��7���_W�p �S;�\���������%��(��L��3��qo�� �vʢ��g����wN�I@Tپ�ڪh�Kt����v��wF~�Ϩ���U���#��+���<^4|O⨣�&�O���V2MD��֐,����q~e(��@�igI{�GTk|t~�\cH&>���A��ӥTG���(q��z�sۃ���(�} ����gu<�R����mö� �*g]��)a�f0*���ƒ����`�6�0�nX{ޚZEMT5�L�Q�YJT�#h��`����{
x~NS��ЍZ�(Q�G&z� �!�!�B6����mx:}E�Nx�l�v{�*�i�0��V�#?��K_3`ki�������	e�P�Yy<�07h�	�%Z�00��ܺe�֛�n��U��ᐏ�
��F���;yd�RN�G�pc��b6�f�3�}�����zw���X�\�X�*o�
�}&���?HdM_�
�q=���a�MXb|{�PB ��6�w�{c OG��������#a��,�R[gcdj!7�@f�)-i��Z2���i��>�������~y���i:!M��VlLxN��V=�b  !��s�A�B�#�̲�?T"ɪb�Z�΅��ԅ�q����u���f�}����Q���~��#�Ѹ�������vE�Bx	��USj��Q�y�z'JS��,�֚[�eTЛA��V�9Z��h~��5���C�^�ň�l}|�]���Q�]\�����W��8D"r�垙M��`���*�i��0ό)SCYX��cĪ�Zdb�f��Y;��e5p"ū���N��y�L�S���g��9��5��>���k���@ͭ9n\��ѡtMQH�� ���u���oЧ.���~��|"��tƶ���<9x=�(��8�q��5�|Ze\��� �e��];�[���n!���X�i
Qk��AS$f<&�a�D���[獑��U<۲iվ������ck�>p���,��XU}�kZ�x�g��ܻ�,��<)�x�{�b0�v����C��w,o�F���]7�=���~��1�"�߭�jS8��ű3���R
��w(N������]�[uF� 'B�
-�x��b&��OO�*(�"M	\x��ȉ��{0��w)<<�<a�\�`/��: �^)?z�>��`;$]�at+�/-5���Ɵ��x�#-�C��ӣ�Q�F�~�b��d�G�K������VɕA�;����c��Q�
�6��g��t˚Ѝ��;h�A�M���P;_����z^Q����?�1Eu- !��L�[�,�wb<=Y�{���K0'@�P�1[�t���???�1U��P
��xE�������ڽűf�O&�:S"�B��p7|��p�S�_̢t ˌ4���%1��߰-+>�����j���7�`<_θ֡�]UϜ%��JwL��[�"�T��'��g�uEQ5Kap}�Dx���w�QC�{�b��-%�!��)��D�}�Hc���'���"���[7(<<�
�r���5j�v�C�-���������P&?b�9�HS^h7�dI�.��D�y|`T�ԟw�^��y�ix4�G�=*��gc�w�$���H&��Z"�.8[�O�~��@���%6�u������:�Q��A)�4e\J�֠�R�ǚ�h5�޾-�#c��HO��^���Θ9^��c,yh}|F��G4�>7�~��bT����$��>��b�S��7�T����of�K��a�hO��������l��o�`�I����3���J�u]�Ղ�oo�]6�N���>�c���)kOPb\�!�<g��YʆRW�ց��2eJ�sv�AZ���O��\�x_߰m7$�%��������% = �Z��L"m8���h��"_7�V��<��~�O�;����˿�?������̭��^ӳ�2yqKjM�D�R����P��B��$��:{�H�����Q�[�a~o�U**�t/���wV������ק2�|w�Ff��1�����|U� g������3B~�(G��{Vܨ >��8�#��4⑎c�c��~��>��b�4��u����h��Ý�Q���8�[�VJ�}��b`.O��8]���6����nn5�f��<Ns�<%�T�T|�<���Tf��-��9�K�����.R�����}�.��\�:�UN�G�n�c{!{�M#��އBx'�Z�H�`�P    IDAT�����h0~����E��8���F9�c��Mr>�u��c=���L��0�y��k<����h��d�������X��b�@7W����e�m�S��#)/�ܐ���6�&��X��h��2�t�P��z�Z�UT��bM�y�vFr��?lVv�DXo7��͠�a�Wɛp)��<�jy���v�y��B���1�Gl�h��0�']���v�g�ׂ��W��	?�����W�o�x�1[���3��|ѵI�� +qIԱ�Mc꙾�Кq�F���H�@ih4�@|�J*���"�>�/,�xf�n����a�q�ٺ�wн�?
��"z�.���edh#��H�=A�ޯ����m�E\�#e���	1٭ogZ�_C���vM���'���7�9&5������Q��W/�
]k֛���8�=#�JǺ�jhV��
ʊ�4!�Z!�u�Q<�	�Yv{>[[�e�!W湡y�������ʐ�(��9�|/��w;{���M��y��?�I��t�KW�43*q�w&޹ϙ:�����g�}`$4��0~v�4����>�g�E���ﶍ�����p�u��1$��G���xT�8]���T�� �j�)u)J8�����V�{|~�àX�)D�t¦��
~:���		d[�P+ѵ;��
�ac(PCtBk�c�HL��_`��i2�ݡ%uc����<�i�ؼ��\I��fdH��{�����o;�LU�����|����<cNg�}{������?�	_��,�7෥/<����
�[j�C��|�����s��y�|>a��!^�#r�Q�U��k�Z�ca뾤δ�������i�-����?Ҷc����,Gk�hmƾ�ew����h��?�ne�]��hA���g{����h���Y�q|�}&�� ���x���c|�ޜGk�h��ϸe%��E�A��u��E��,�������v�����V ��"�!�t���RV,�w��!1C��ۺ`�O)c���`k�<a+R��&�lbR���������-0���?h6����1��W���߯�sLtP�
Y�51$�F%��4������3���<�O���<�]�r(?m��0*������U��a8$�q0>�y�V;t�x��}k1�gr�V��f=rx�=OA��yϧ����������!"ޞ��<�m3\
?�O�_noXU���������Ox���9!gC�3�8��u�D�mYfW��H�%��PIk'�Ći\�bMb=[x@^�	��g3Ζ����\�ND&�l�X���d:.�}:��4���M:�}���/���?������������gLH��j�Rp��i�!UA��IQ���9[B�X���j�r>�����&�ю�,��R��`#p�)'�)l0�U��Ǔ���u��>�eV�xzz�z���3Ax�Vp����A�%��_�0���=O6�<k�w|F�K����"g=�-?0J���ZGAwdlq�b��H #˲�F0� u��a�����LR� o�6B��e杠�1F�'M{��;FPz�o���E	�y� ���iw���9��n�RBk
B��/A*��ͳ�m0%��*�u][&x[#�5u����
�UQn&�O���m{���}��i��n(�����Ԃ�vBUkg\��2������yB%�LV�^����e-x��=�Ɏ���S2/HRO��v�m�pK�#��
)�LJ�]kԑ��ڳf��xX)֟;���-G�^��l�2�\��Ͽ[l���Z���7�Y"˅X���+)�^�4Z[��6�b��0r�w�}��AT�ڀÌ-$nVx���(ۆm����5=��uHK)a�g+��C#���*O���D�ݶ2?!�˝��V��(�s��E��!>N�	˲���'�%���ն7A͖��Е�JV�;3���eG�ڤ�~����$���Ys�H��ॼB�����T����o�@�7�TLd�"��^�T<�����u[��f��)g,}���h��Fa/�n�O9AQA�pEǺoB_;�z�ﮝ�G ���M9�|>cY����p��ϟ� E�n�����f��a-g�\-O ���HQ<Y#x]7\��ۢ���u��BJ�H{W���{w�ҝ �����k�X���?���Ԅ���>G�8�7���b���ނ�4A��i[ND���M靠$��4aLC��zŽ/��X�#�8J��K��	�!Gdt�?���ŗ{��w��>�Y�6ڹ-G�M�rPF�kL����ya�6����5aW\E�b�����"��f�~�8�Zb����f��e(X�#�}��'�%��
)��EP��@V�>0J�Ԋ{yǧ/�AS����R^����b�Nx����\]Q�΄Uf$� ����ȧ�@�Ȝ Jr>8��5��	&䁞2'l��F�� VX$� �!�-,gۧL��	��!AÂ��k�L>NA%A�0'/x�%��e �h���ֵy��}p�u	���4Ё[�s��9#'�xS%��x[r��g`ʉ�᩵���E��J/	32R:{x��(��ɀ�R%�r�Faq�E0s�iNͫ,���mk�����C8���TՔ����u�����k�(J�`������^n�x,,���f�\_�lmKmH���������S>!c��DJۏ�S�������xH�C�=[�l� "1N�|����z@s�E<@a^�'}p=t����i�X���� �w��Y������c���7,�E+N�8M3n��t(�SS� I�,�LU�n�g�xK�X�❂�I��ԑ�
v����bN����b�z�v��Ȳ�K)X���>
�х�RO�0B�z*�`VH/�	?l	Wm^&C�u�F%��W�P[��0�IM+�^��Ƚ�4�[h(�|��/A���&ߗp�h�ԑիĻύ���zp��� RG�:
z"��废��8���NA��=4��
M�v�����$�?⟪YǵHc޵V��C��*����ļr9Y"����	uٰ-��"1�E5Y���6�	�R���/���O߰Vã��|�9M(ۆ�����;�Y��}�Ή�MO��nb�lu��Y����XTRQd���iF�7�!�4O����o�d�T�rr%���6He�`�]�{E[>��{6���A��m�ߟ�����^�X�򯯦��Ihʬ۩u�r�MF@Y���������p�K)E/��b�W���9�Qk�K�r���Y�Wj�@klD�[�3#�w���0�"1'i8�4e�4�{~5�~>�����ij�6N[1o�&k�j��B�6\�E�3�Ɇ"�IM�� ,���9JO�x��#e4тW���UVXٽ%�4͘g�v^|��b��(�{|� Ӓ�b_�}��8��+S"#��≞�����Vp}{��@>_���_��������S���
@;]���X�������3f�o(7���|�`�w¹[�V50�5M�tμcr����.^�Oi�Cv�>�!��C��	Y��{�D�z0��U�P��<!�u[��7s�eƩV\г��G�|���P�ink:��=�Հ�I_�P���S���`�P$�ܗ����1��Ϣ�����\��oއ �	���y�{���_b���y'�F���eF$����bJ�5)�䥜3ʺ�v�",GF����ܦ)1>�`�V�ui�yf��ҹ!�?����"^��������?�_�|A҂o?�����/�~mΞ\Kd����;F'�c�`�����#|�Z��ѭ,��ɘ��i&OXTq�C���3ji�22��Г�Hݣ'��U���D�5��V7��z`��֝��Tr4����c�g*���G��:0�z����EX,�\���c�B��˚�(˭�L5O�AªZ������c�wE����VC�'u��9`��%Vm�P�:}�g7��|N���g�P�6df�\�P�%o� Qv� 0o���`����˚�Z��U��eY1A[�<t�	�<��=�S�1�qDR����� 
������=����^?�d�*����pdq�\��nՁ ��vC�&�s�*���;��'Pf\>¶mx��7��yrT!�� ���o�j,Cۂ+.�>�������?)Y�`���o��"p׮
ΐ��
a�6O����#30�cE���m�,��;&�PE���œ[mJ�$ �����e �i2W�3i�m}��\��@*����Ŝ	�DH)#q�1Im��
��˚G��Iw�63�Xs���d��COw�5i�E�(�Lk�P=����Yo�	$���i����۠o���`��FL��3�N5��Udv�7fT!L';�y��3н� [W8Ƶ-�`>� �I����D�U-�9�R�IP�qb`�����1X*خW�X�Y����T�>'�P'լحVc����L��yƧ����ח߰�����NV����L�@��G����]n˨P��x�(�x�{KvEW2�-�t:�gh��]8G����.3�S��}M�RU��)SihDd X&<7�+/􀡏9�X���';�?�A��u �����ORO�K�J 7�^J�-���`��i�sac�gC��m��@�����A��B��p�!�2�X9M����njFv���<���"<��i���/ϗ	��	˺zn�y j
�+��\q(-_@T1qF:��nX�Z��l�s:M��`������"�M�%�)����¿{m����㪊�2D�2(�XI�m�jX������oĽ���V�;���ų4r`�wS��z�{���;n�H�쵺�_���9���g|���nx_�/}��0�8�j�H�Sǣ&2��!���]�/�u�^�Mh$�j~��r��h����~/�zŝ6mkʃٻ��D�6�v�wt�փ�e�P��(���!�����,��K�]�i�S�"I��UP��9 �ʌM���!�ld�m<"ؖ��Ƌ��.�12�+Ӑ�'^7.�����Q ĺMя��`�99�6�G��h���&ޟ�	�u�O@�R�׷7l���!��_� (��1#���Ko �D��B�Z�e��ar���n3۔&�T���\���lf���PϠ�%{��)
&�RŴ]���oo� �<B�����ځ2!���!B�h���V�ؘ��ܹR���2���k �h_�Aǔ��]wk���81EM���uxE*(BC������emkAq�$P��@u�0Xڑ��!Z!�=ᣄ�*�*��C��2O4#�����r�U���ĂD�`�3�Z�:1�����f" Gba�2�2�D pRL�;)%�zgv%���<�J�{(���w�uzL���~�Q7z�JK����ё[�)%�9��b�6ɺ*Z���z��<�[R�T��y81�0�&\.Դ�v��������4�p_�%ԫ���,G�]�Τ��<�O8��r��ʾ!���\@s�������9�MG&t��>�r�e1ANF�ۺ@����w�������oXD�7װ85�$C8U�O�g�{i�� Y{���)���~?8�N�/z7W�\;���D$W�$�Śk�?Ce/prT��`�r��b(���.��:"�_�:nڳ<����p�!�L�A�8��͘�GVғ��)T' �s?١��V���V�#o��S|�<(|O_`^�O�Ǔ���v�Sl-�}�ǜ뺵ܔ�e�w����ucm�,��SO��	Ĭ�/��v�,��� ��^i&o=9�a��="Q�܍k^���!$��)c��&.b��L	��@�*���^�9e�U���@���[�~@'c�|��0)��W�l�D�X�(;�F��*=��-3�4,���+��bw�I�n�@���Q�Y�F�^�Ϟ�K�aYq$Q1C6��@Gae	�Q��^�6���1D���F	��⥑���\4E���SS²����*�����)y�&�ߦ	e������Q�)SlB��#GB)�Z��	�}<& ��ɒ��R!>~��'�ӡ���I��F�:v+�Xk1m����mXw߷ZQ��JE]m�k̿8̒(�l��r/c�օN3!Ô�$ /�
>��kԔ>����L
�8�(�o6/�yS<��t���G<��G�O*A�La�f�߿zӐ�]��|g�J�8�NP���y�0M=�\�䄷�7�����H���+�B�Y)��QC����41��������-T�o0�����4�D�������Y� LH(��E5���Rs�޺�eu�>A�P��B�\cY���W=ɠD�H0~����.��ˀ�!���C�20�YU�P�ncd"'p�R�V�8h�n��t�՘2���` �Ѷ�m��h�ʁxOf��ehS�`��a �
h�u�>�;/�h��������u�Ҕ
���=��x4V�YԤ��&�[��%�A
ST7�>�jD�!n���E�sB����٬�)�ml[�	y�$����E?�J�L9K�Q(Œ��c��y�|��m�ۺ�}V�������|��dess����j� ��^x2��`��Z-���Y��!5E�x��B	��{Ќg�bU	
�PJdp�:���aoE�c�����2Z�$=�
UkD%�\��N���6E���@ ʖ'P+R��m$��)e�D���|�+�d�c%L��
���w�S����]�*�Tf�
)5# ��l����
FBN�4���o����!��&��RB���W/;~��qUKЌRC�!�2�C���y�����;� FN�ǵULjr�� �gLj�Jau�&�SJȓ��H��ٍ��j5��`�[����PC���nmq��:-АU	 qM3h:A�����
� /[Ŭ�R6�s��'"n1����O�H.ك��`���ϔR�?ew��k/9�i2"�������?�\>������?�����?�T����,�y�l��5;�����gs��% �[�L��eG�'���ws4�!���
��yR :�)�[ת:�<A��i�c.���R�JP0�j17�L	k�sxM��4
T��+9��!Զ�꜆29�ņZ�����豤����a�wU���`ϥ	U��*��%;��V�B(�������6GN#@���G�[��h h�֝�w��.!�=�,��� ��۴k��y.! �@4���W�Z�s������A	L�+�l)��u�����g��ī;0B�8�8�@m�����3H2Hk���)��;ݔ����.l�W��^+	�:�\*�zÏ�7���!�����Ni«�������Sμ?wN@�f�[\~�{�_��� 	U-DݲB6����Pyq�+�� ���a�Lp�p���~���r�%��	�c(��x�^AG <��s]�e��/c&Ʀ�	@�Y���<������Ah8y��w9�(c7��1��2&FW��#��Ϙ+K�	�2�*
��p��\[��E#i��M6�@W��[BS&��.��DZ�a!`�V�M��C����窊�2�1�UQ�"͌|�����P�(��ʧ��Q�TKf���3<�p\0V��0������>ˊ�ނ��N���x��������k:#3��l6	r���}`�j��=U��f? <T���>��F���VWj%)�
טZF��7�*>�(���׭bN3.!(��|q�:�ع~wl`��`�-�6�|�]�މh?K�=Ӳi���ۧi��8�iI.g�kq�)\	�^um��A����1|b��H���Yd�H���i������eI��j8�+H��F���&�Y�/��@��lZ�֧I�1x	�4�؜���c�Bڅd�MN{��W0�8� ��~	�L�BbMQ���EC���1��(þ:�*5�a�\�&`���<"��Oc��D�3F�Vcp�E�$ȉqr���N�%+���P�~]��x?��9�lm%<<�Y���4�8CH���1<Qt�;��Q��Ky\_�FK�N��xT��HKV�~W����x�z�^ۃ��v椏G�1�}���C��@a�ژ��L��Y����:9����3
�=�6�6$P�z,Dܚ\F��  �IDAT- �E({5�B�h���0��K�uf�wY%"��a �ʦ�	&�l���,����7K>��\T��@@�9C��3?�A��΂挚�5l[�) �\�e7P�
�'!h2�p����Qx���_ΓR��#�<6�J��-O�����u�pd܍��Dd��]�s�ܠN�6:0�n-v��Ta֯=�]c��}]��T�~�g<�E���WR\҄T��<>�c	�	{ws���@'l��+���R#'���� ��
j���dnF�1jB�q(Z��^y9��Q��jl�B͙8��XN8�Ćy��2�^i���wc˺+�(h3h���7K@1�>4�ZA ��u5��nN�>��7�X�f���n!k;�A8w�7���L�J�Ad9�:��DDK����v�Ib|�"�^51l�{�ks�z4L��p�P e�"��c�*$�x<OV�TE<.Z�<���B8	���i��ۊ����g�цӔ�]V��
|�zd<:%sG�C�4���c�1?�����)�q�}��b�Ċ9�/�p�#��U�;��Gz<��68���ϴm�\�=_�g(�Pt��iw��M�VA�<]�P���x�"�5��Ce����^�Q�Ru�k�p�>�"'\T��F�S�6�2a�d�DX6���ЧW*\��X{e���w���JQ(�ܕ��7g�Q���j��;���6�ו5g"��z�L�7Ο��:�;SF�'���n=��c�U7˛"Af���@V!(��$�����h��ᆌs�1���׾y{"r��ܭ(����Z��C\�dI�(*~���4czzƪ��톥n8��7l��	���Hz�E�\�Q��V�}��l.��0�\m�ĀE,��ȁ�T�QE�[�l�{co�����k|�6�Bu&�;暧=���9YC�wa2��Y:s�-'��?&-����Wv�ʐ�2�gk{)�0����� я=��`��X��hBޘ�P/M��`ަ֖��
D�)��.zDfL�{v�p��ؕ[���.�ݸU�i�hW�y�[~Gܓ��uM��f S6����LUI�q�m�U*�j^*���-�$�
Xo�ӄ���Qkqk���,A�֣�M,@(��y�Ϡ?ZS��0�χ}��l��fl[hw�P4��H�w��sC�+ ����~�tT��5d��P0R���Rx>Bq=��<y�Wc.K4=8?$��W�1o^/m�.(Z�,n��0��ڞ�#�A�+*NdȂ�<#V�&(Ȝ��䲊�2��z�0k�0,Y~A<[]ЗemF_���&T����H��0`r��`�9����F��ذ���4A��`��	R7H��L"ji(�-��5f�����!�9�z�߸I{"���Li �������� �+�9�Tv.t`1	*
�
4%|��>��=^^_��_�"XK�n�CJ"{H �}�QB��˔��1�>��=�M��*��%���Q"����6\����N��;�(������]3������3���@�[2Ҁ�&����rʸƑ�N�$���2�4���ܫ��R�
�q�C��~���qӏNׇ�$�u'�&�,I�JkH�b�.4[y�0�ȄQ�q��F"���9m��9�Tq���)��\��X3 ū�~���1%hN&�iF �YY����
���
-��A������5k0~�;��"ޯ�6X��G|'�gJ?R� ����v>�TuX�v�DH�cgG:���Y)�*������L��?��+ ��ǽr��ų�O�=��I�����a쨅q��=0�qf���ĵ���{�ΘXED��&��ھ��}�����-}� ����s�1ި>�u~��Y����(afF���	P6ܨ4���H�� �������z����c{�]�W���V��e�<��U�l�b�+V�Pd>�@�[ʘ"{�454�m�����[3�Ljw���[ܶ����'# QGs��+ޯ���໯����	x:�T�-k�4=����\E�Q+��Y��K V��ś노�.Vs��У�=���	A5�mt�vd$�����k�nws�\ss�&�C�-#<�=E���h �����9�&?���P�/"��� 3�i����.�s�
�4{͕*�q|T�0��j��;>C��cHH���}n?
́�f���IDݺn�����\�Z�*j9��{5�pO:g<}�����/Plxbë'b��L9NS�v��(K�d���9��{�.����u��b���u	��Ev�< ��OӾ���'v
ذ�ad�r�hWx���>���t����۹�n��(��d��GA_x��x_��ᑈ��M顴6�'��=q�!`��t��"����sl�Ͼ�١}k�(d�p�	��n��`��g�	x�\��c�F��$�i�M�*�g��qef��*��8L�  iI��� �����X>�������=2M .�(cN�@��3�����'��mJ��n90�A�v��dD�fY�J=>c�O�e� ���6�	_2��`����}k� ��N��/Ӫ��$�1�f�:���D��A]D����%^�<�(��ql@C�S���8\���������;�E�����VT�8DP���1 �R�al#S���Å��PWϦ�A-㨉vs��XYN0Y�\�1��c��s͏�zI�=�[jX�Q(Ž3��\��cc׿�ʎ[luPI-�����&��^�cډ�\���J��Yם3���	q�<��,���2_�������?�_ޯ������G��O�'�<Y5��DK�#�z��q�Ci�є�(3�<���r|�z�@�1���=�{�0�ȃFC�d�I�Ù�>wf�Ze7�ݝ��S��$����#�	 0�5�L�*X����}�����#�{�)����{�!��\X,=u%B��O;�����L/	�jJ���0O�5VU�K���^�j-ho7loW�Z�$��j8%x���`j%ù¿"��7��x�CV)Y�H1�B$�)�^=P6AEE�,��A�Į�L�������K0Q(D�3;ǣn�_�Fh�C�Ӟ��B(��YЊ:�4
Ҵs�Mq9�1C���Z�j�i�P���m�g���5z��Ǔ���!r�-`GJ�R@z��#3*n�gbP"Is�W)�A�	4~�@#s{E����%Jݟ��v����!֕��P9n��QA���ZV���F޾��X��S~ڽP"��#�8�9 �:����|ݕ��~���d�"j�T��=M��&�����:Fj�p+}�g9�����!
,rS0����ܔ���������:�6�P�򽗩t��wBr�gC>��'�$FD�d��[�XP=�GD��brl����z������[�?�	�|�kz����� oj-X�#��y�BЗ2x<�c�7A�����o���C3�{a+moƫg��9�%2��@8*Kap�WP�s��(v�a.q���b���ݹ� � x��p�Op�I�ץ��p��0�Ճ��	����k�
f���X��ⵧ�l��7)^���Ҽ:���Y4���t8gcg<���u��&<�Y7�{0^&PT�P�BL���@a�)f;k^��gD�.�Q�OɈU���31&N�(�����������4mr�&    IEND�B`�PK   �x�V6�0{ { /   images/c51b28eb-c857-4ce7-b81a-d633a3d7e747.png L@���PNG

   IHDR  �     �PVo    IDATx�	�,I]�U�U��Ww�~Ι��>�̰�* 0��p�EAQ�^��z��}W}>?��wԋ(>D},*��� ���s����]{eVVf���#�������90H�铕���A`<n��ݰ:�t�������꣜�=�3s����VG}~I��ԗ���_����X�K����e������{m�2lA��"��(�B<��rFL���8"A(d����B�"�R>�
	{����b�o��xݍ.t��Y���������2[*�E~���$�))K���ߑ��߷�[7��Q�CFa��&�(�[{�dD�\{��K_Ku��#k���d�d��^�u�ԥ��:B�>�+ʺ��L�R<q��蒆u���7ц4ѥ;R�]��ߑ�t_��G���\�HQi�8~��P�z�{/����ne�^�����S���~�tA�y7�W8Nz�f�У=u�Kt����j���T�%=R&�9��ߑЃs�8��hq��2.|��C�n�?yL���<^�/�׽F������+u��2u�[�v��d%
WA�Ks\W�n	��_!��Z�N����>n���Xle�lu�z ���E��{��jr�"��+쵇.ȻT�v�+*W_�F;$G������(�:��b��vC�'�����l+�ӻ�xb�a;����m�NФ�<�@�ʻT��P8���o���>���0�z�E3�\Ԍ�v����p���g	B��(!5]�q]^�i�M���iEt�����"�G?��F�P0���A�k{���Z>�g���-W����O�9U[_��՚���=��[isշ��7��n���J	��P�,���ns��b1�I �0�u�
5Mb�a���V�"��F"fh�������f5E	b
\�Z-!ON��\Rx���&D�F�Je� C�p*�������}�{����X4����xڊY�*��vHU��~��«��	?0�$5Bi+dm(��ԕxk`��I���Ӫ�_h�:ҬSRlO��M�IZ)^�+m�dsItL�j
|�A�Cㆽh��}�%�1����u��������ז~������a"�58'X��!3��~��'&Ǯ����H��+���W�,��BJ�Ѩ.o���/7/���]�n��x��G���?|�Kw~�q���d2�ڑj��(��f��9�_n	"� {���I 3cd��$�������-��\,b�[��3��z�u &����h�uG�{C�N���O�K#�E�:H'']У ��L��Zl�E[{�I�Zw���������'-0l\��C`*0��:@QG/b��t�v��9	�N]�^��1I� 4=7K9r&j�by����u�P���a��A$yjt��sa�d�r���H�������?qq��6����ly^�n׼�cG �� `�Հ:��P�"��n���FŌD� &E�F�����i3�m��@w�@�n�à� zӧ<��{T������Z��=����>Q0�D�3�[|"i��o����=��F¥tl>����P���hD�h��Rw�A�x���^���c,3��線`L�5Ȗׂ�X�߼���#��k��� �P/�!�4"���:���Ѳ��g|����_����g6� ��Mp*��k~:��g3)�S���Nӫ��57��B2�����x����ut�n�7���fe!�M�tz�o��]��A��xP<䰎�^	��61���P��M���������'� �#����V���L�O��vgkp�JR�<-V<"�0�mb��l����1����f!м�E���6h���F����M��~4��v.o�t�5@@)2�V�@�^.A�h�����w~�G�~��^��M���v��-+X4]�K��8
�"m�hS+���\vă�l{��,X���R���0�i`b"#fG�E�u ��hLx���6G3,�[�v�H����ޭa���Ԧ0T4�)����`�l�c���;���;V�-�xp��r6���7���� ��8kr�LA�lk�#=�i��
C�d��#�09aR��O�L節++++�Z��w�5::r���M��hYV?A�S��������|�����B�0�G>��;� �L:΢dah���"7o�2�|a+���cɈi�맵$�ZJ:���Ax��pgCy�]��ݦ=�a��"юt�O�W�p��'�e�O��!\a�,�ȡp�<��z͵������]s	'g;<^l�}°��ֵ�H")���8N����¹D�mD�_
�X�p,Kg��z���T�V[��o\y��7?}��]��{#����/g%}��[���گ��W�vw�^)6�2�La|�v�T2��N�C�d��������\��'xn��D.�ɏ%YGnd��V����2x���*�08�/}�����#��d��aF����s�R7�j�Ρ���'����wPZ�F��>�ȓ*~���������*�����W�K\"�Vm!�,o՚���p#��L�x $��:��6\^^^]]-����8�w�0���d6W�	(�|&;5Y�֗=ro�.^�k���+7�x���H�٤���钢Yi��9B�9����l��x�\v��-�^.��3�'��ؘ1��,�E�d�rzeuqa�t˨D�Љ�a6��A?�C�j;v�aׂ�s�Lv�����t&�f1j��W��휸�+6(��4Q֡!�_ݬ��+����Rj�xE�Z)˶�H<ƭz�	�Q�i�� $���S���5'��P�����36�$��+��ģ[*�����>G�@���Af%�R��4%��|�h� o"MX�="M^6D�hs�:m�50f���V����#�����ﻦ�}e�>��6Mj�cs>��H�Va�&S�Y�Z�F̑l�ݮNF[n���{�����t�Q��n+7۶���[K��'�g[�x6aeWc�h�����_ر���J����ܳ����y#���v�������T�J%�c���5�ż�A^�;�TP�Ї>q��ii��Z-(��hԛ�T:7C~�Z�?}�a4sik���hjt,7�{j6�����y�UGg�Б���B�'��ȏN�V&�!�a����BvT�Ff�5D���.Q�?��p�p�.bCm&�h�B~�hذ~�0�����# r�Wh��|�]�e���#U� P������@V���2�31��"e����+=e�5��)?�H�B~R=�}�n���P�Ѐ��K�i'q��m/��@�8e��q��u*�'�:$N�ʫ�]q�~�ˏdS)��ٶ�!�N=1K.�} je\/\,�V��MNx�yͫ����ۿo�m����x���2���e�G�BMY�	�4$=~|�c��+_Č% =�P&���@n{�y���*���������7���!7�t=�)[�ɦR����}�|��嫷���rqծUw��K��w<ٌ� �x�n,�����
����' (1H�C�>) ��B6:�R��D)���v���L����*��te�uZ�C1rWޘ�V�TB-�Z���)@}� �e������x�s�����-p�`0�H��y��",y"A<;v��fm��w������׿�U3��z$-�t	-O`�T��J�������?2wf�أ����+��1s�Á�p�O|���������"3� �erQ�:'�e G~�7��؂S"�v}�#��V>����?���&&'�`&���j��i��|.b����w��^��/�ǐ����O%d��e�M̏�jzj�)�?�܏=^�V��X6��H�"�CDDwR�R�)�R^�DA�n2���R���(�l�L3iAf�aH(Ey�����&7�(���4�y=j�����!�#3�:Ga�L@x[&9YqHX��IE�q+I���IR�B�nk4�r�5�D�?X2.���v|����!Ah)9u��ض���d<����9���n��w��������4��t&���d90ڳ���x�E/zn&����G�%�j���B�������4�Lv��� � E���V��]�T�Í �r�X4~�|��� 㹕���,�İ(h'��F}y��c^`��/�����/�r�u�(T�B��rAH���r��!@�h�g�r�����3g�?\�ۙL:�����͒���c%�R��`E����+"�9�)]�6�t�%�9�JY�d�X�@��VE�H�m�������?�L�@/���6��H�`�r�t�>�54F���}LhK��-KZ��R+)�h٪��U���خ�vl�ap	(�k�$��f�V��2��|zuy�����Л������_}ֳ�g�>Xz��+<H� ��fӍǢW_}��W_�R*?rdyn>��
�w_x��GW�Wn��i�Y�i��mtQe��������l�\~
�3��?��'f3����k~Fk"V�,���ܩǀ��������V���r&�H�P{"��2
���?��'X����_=9=��~�?�9~v�|�����"��
�\�'��Mv1����S�M��&"�� >�nԝvPq+zf<�,�9齥��$����h�Q�8b4�s*r��:��� ������4`���,zDV�ދ�>�n���P0���8� `��H�R�=}���[~��~�W߾o�y4l��,��Q��2��V�r	y/������v�׿�/.-�ݷw��@t=֨��q����{��et,�#t[�l<+���W�A:��E_������G��1BV6;i%� qs�,o]�&��l�[�g��?�J��Rej��˕b$J%R��#lа��)0
�{��je�0��>�W~�?��������Ri<���$!�e!��2yv-h��k%�Y����m���&4�axí�_��F��[o��kީ���:i��P�Q������g#�P��b4��D��>"�6�F�`�Щ%���惯�nl�[�{�zd�EV�C�Z��a#�J-��5ȷ���x�k^V��J�2#\Z-�G3����x!�D�`���1��N9�\s�����?
�v�w�\vM"�Md'PO�ҝ_߻o��_�B�����%�q�@�(n�N�������_�vw�E�0�2��4��)b��~ear��?��XL WI�n�z�Dr��\�P�
0�l�1���|n~��������O��/��]^�/L�J������4&?DY���h��V��a����Ukۮ[m������˱S���=���#Ҧ��+j��H�L�NĠ
ȃB�q횈T*�6aZ�_�2�@Q��4k�2�]m�m���XtF�E�\b�"Q�����"a��W���~g�e��l�4�{����bI(2�8t�԰�#��"��{�������q��C�r��+�������c����{��/��禓|�a1���4��+���?��j=<1�/��,�	��ťs�,�A@C�e��^F�z <�	"bp���ZA���� �s�===�a'D~�~�СS���ʞ�T�X,F����IP�:�Q�򼮺Q_T��(T�)�b��8N}e�bE��g��� b��ُ*�<O�b�C��'D'�����	t��d��LDk�]CP�-���r��b ���,�C�x�Ş�/�K��GϚ�1��Z�D�^��ZZ\��۽���w�����j{Z���A%�]��u�vff��++�	�:ƻ������;�E�Y�Ht7@��e�`9O�8�*����}�{��u���]-aB�L�:�4WVε��_��7n}�7�@��%��Z����;�e�Q��V�4�oTʕ��#��׿�'����D�����\��T'�h��ND���D�ZNgR���IZ�x��?��/9U�i6�'hCR⠩���~T� �׬�8y$b4߄v��_��4�������� �~�"+���6]Xb`u25Ѷ�� ]V�DJ�/F�BFi�6z�����~�_o���$b�����r�'X��w��>l��v\D����{qi�m�Qn~�����=S�R��U`?ht�B�^�B� _�uj*�<���ר���A��G4�Ņ��y�G��k������@g3V.�T�ъ	7�V��D>j�I�RįO���{���?��[�5:��+�d��?����ALUu !���jd�����\���#G��
���L,��n������Z����E��n.7��ڳ^1�z)71�]?9!���������D�^ k5b�#�s����W�XDR`�מ���V��;P��R���#�Q�r����ӧ�V���v���$��=��jq�0��L!�hH����/&�T-#'�a��[��-�0 ��]n7�b��c��[��������~d`di��?JN ɣR)R(������l��NE_��������ǖ��kK���m�̙s�S�up����/��d*Ui��
�مw�����k�����=��d�!0��I�\��Rn��ĳ��<V��|�3�����2�^nAW�ڭ���.���GLu�KЙLJ���F�N�޷g�e���������+���M�M�Y�<��X��\�?s�y*nœ`$�-cm!�+�/\m����G�P~��)ױ�����|���>������F�F:m<��7|bfze���KyH]ժ�Dw�S�ۇ��n�-� N��mpU���ܽg��/y�����  ��R7R{����of+H�(۶19}��_{v�g)W��S��X����N�z�?c�4���$D������Z]���1tVKe�DãH{�]�lJY�
$D����V`�EL�iZ�80�o�����#(@}��@K87�N��bC���5�4�N�(.' \�Īa���,ޙ�qߙ�}�{�+�p2�/L��i$-�N]\\4�P
�<ZH��9]�\ȷ��r�,��V�����࣮�X��կ�s��3�Ϻa���^�7�M/�.B(ӀǦ\RW�`;l��v|�-�g	��Y�)��v.�,4�hd 4|������4��EOX��G��0Xs��6��Ͽ�>��3���ꃦ���D�������_GF�VΡ\��0�~(���l5ab؂�5~�0��ھ�DE>�F#J	�D��<J�Y7I�r�sEg���������]S��$��k�E�2ȗ�p����p�=ҍb������m�өĢj4D���['��=}��H��$�u����f�i���I����S+��ü��#L���D&����r�:{�\uu1��y���~��u2�*�v���9���H�D�#
R�%�	��o�r�.�M��0�%~�h�P�O��e��P�5�!$I4Jj��6|6_TtLӌ�r9�g����RX�(�o!�x���-,��C�������Q e�\C@!I���Z�|[��8K���_�kL�e��ѻz��:�z��+9�5EшT���LNl��h��_�V�qh�u�̓f@u����df�� {Q���3	#��z,i�\�=�p��_ͨ˾@�f�v�
6�t��]��>=pK+'�d��1}W��v�uc&?�ctlO25u�}�>���a4T��}���P��d��V:�dne��D�"R)*��" ��.9|�a��[��Z �c������p�Hi��R�"��/ �0R�g���$�F!�'�Z����7f,�����h��Y��Ђ�����֝��L!���	u�3��N;Q�GQF�D�!N+ڨ��JE^�%�� HG`b�tꐾk���.hv�b��z�T5��#�w�Tcx(�;�r(\j|���%���D8�W��n������ફ��Y\^f$Ԛ
c9�K6�:;�
���o����>�j�..�M���^k�	�����v�O\ML����{��ԙ���|�^i՛��Uh�dr�/Q*=/��j�R	;�&����`8�V�ݒn�n��v\l`����X�!��ë7�lRi���P ��Q�&wb�ۉ`0ZQ��-v�d��[C���\(;� y�p^&��2`��*4Ӳf����6��8���F��    IDATx6::��xٞ=+sgw�G���𱳪`a�!O��!RE�D[<J��-+U�S"a+�H#7MXf+ix�����I+������W2Y4]ن>r���)�����T�\w��5	sE�����GB����ڹ��JdR�V����F�jz�b��:����S_OZm�RkBZ��.�.#�f$V�L璓:�����f|��c��T�z�������U�<�g�U�Ӵ���E�;
��ʹi|[hZ
�V��V���#����Թ��۪zVSJ���+^џ���k.�:i;_M_m*>M�Ng꒾�w��ټD��,��%�P��Ň�(�����b�ڒUu}��[�[w�&����9 ���|-ЬV�8�{n��.�I�,.����"�������z��Bp!@��'pR+:2;��Ul8��k2��j��2J�4���i�qǮ>"|f���Oҙ��QH7��Kg�x"'&� *ӹ�Zy�m.X]VJ�Ȉ<h7�b��
VR�!tT(��.stfz,�E�y�Ch���k�"��%��I�h��������! N3��hOà$<I�m\���a�bW9|�:1�G�_��f{������X<?���HQ�8m+V�&�.A��͆h�.JH����Vm�4)<��P�F�
n@��]N�[��~/[{���V*�Q���[
�OtQG��..��.(KV2<־�~��Oc��Tk;��p�,�ڨc�]L&��Y%�ƨZ,��J��S�l6�#3:�P��=U�@�峭��,iqhyZ�F��lm	>�c���j����ۂ?
B^�����4|���ÇW�/�ĉd4�4&)y�T�ۙƹ!��hG�&��Ō�_��m���{���م�5ޥ�V<��N�1�+%���S�Q��HK$�o�k4�-qD��v݁I�Cv��(	�*�N �q٨2��޵ǴB1c	y���e��Vv|tb$�O���NzN��+���-� X����U�#��	����/����ˉ;��G�P:���	u3���]�U)TR�^�q:}7�p�U��!'��V�~�Yj�X9\�o'S��+c~����
��YSѪd�+�t���!w�u6E
w���!e��4��O�KZ ���b�N� ���Ż�z��]�2v��zlt��X��!��\����Y�^苸id�ð��O����9f�P�!~'d�j��<�R�T^"���ղ=59^�ԓ��Ǐ��{����ί�.�K�N[��ZMv�R���J�8��TN����(�yP��Fc0.��A��S�f1K �������Ga	�:�G.$HY���I�F�(u&���7��$LDc�t�<�t&:R��s3;F=���Ԏ�di���}�0�A�(l�֤��6��~�M��g}����@�Y)-3��ڽ�f�
�&�m�`�TD�-u�WW���D7$��\>�ѭ�t�ԧ���A��2�뢎(#�&�8��
%e6�L���k�̈́��y�֗�G�tzϦ���Mq�߾@��T�n��{{%��������]L�Ox�J�o�"j7�^y�{(8�R���=G>���7B3��Hfd5u��G�C�7\��^�P�F:&X	����&��|6ިο���}?���7�
� 4�bdF�`��GU�'��½J*rt�0�G�����!\YΛf���W�NV}?�Y�f\R�g򒱤�䥴�F�n؄��اc��y^��F��� O''�ʭ,..�����D.�t��P�Ie���p6g>t�[G��1�[�̠�:�dvT|Ӻ�2���l�J/����ʭ^���C:���N�ݻrGǮ���J �-���<�	27�Φ~��.�ϲ� �]%�/�	�^]8ۘ޵���{R�n�����Z!Uʵ���O��-�bO�&>hٞ�hWW�}����~�ފth��z"!�`ܢ�}O}���D+P�;5��H����}�C�a��d:�ʲ*�}9��w�5����피W�I�K+��Uʋ��H������?�3oHGs8͵�ڞ2�۞SwR����ҕ��۬n��z./X����z���5��x��	cQ�qXY�_Te�Ee�K����D��j��%��G�=Z/b��ˋދ�F$p��j��������_K&�s��={�\\���Wy��v^s�S���3w|��w?XZ)*�#D{P,�}�_���@_I<��?�(�+�D'eS�Q
���z����vk����/�>�V���jҺ��H{�5T���*b[������P$)���ʧV�6P�.�x;������HO&�&v�-�������^����ޝ�[2jY�	�͇o�+�J�cg�u�t*I��������#)�ht-pJ�y��9���Rl@L��4��ln���S�ڱ�'��W�����x>�ȪQ!�Ej��nO֥��.PJo�	P�Lr�O}��?z�`e"791c����G�0nU4�m.��(���D���kĔi����\��3��v[e�Y5B�J��u�2w3=�E�t��V��Ri�\^(W�q��#�#�p]�kh��#�.OL=|��1������]'�bN�RGO3ڶ=}��B���NQ�[wƄ�&�ꖂQ��[i�u����ڙ��n���MO��y�3����/����\�A��$��������<���RY��	�/��/�NP� WO6]���z��AK���J�:4�b����Tg'醟^��O6�l_~;[��1��M ;�YV��K�`������o��W]w�^6��� 7Lh	k��UP>����0N�a�������:ۏ����0jO�&T��u>�Fu/���!4B�K:.��-Ektl����o�����}������:�|,���T�B���Ĳ���5O�-����S�O��<Xo4�Og��tVzo��=thF+c�F��p:B�c�ݮ���`��0�8����+�x
˝���z#��_#�����D�1���WV�W1rB�8���]���{�[qi��1���$=A)�P���w����d4��dߩ�{�z���|W1h�s(�����sdӤ�������x�Gi��l��68>�������؉c'��,��,T*-#�����>���+�G����DcA��w�'H�B<v|���_:����'r��e�ؐ�kd��]?��-9��PO�C�63��QV�ۮW#fRx�a�w +˳o�?�+���g^]%�M�uY�s��Qtr��������?�����0A���,�ʬ�VQ呢�q�#]:B�7 @?
?L�@M"�����ryrj��N�;�ODC�8�4�F���x�����c#��&rll̲�!���^-,�T�}|�|pL<���;�y�M��'�Iӊ��H:�YXX�����{�����H�2��dM`�kZ�#���{"`C�����P�"z ���Ά���I��<ZP����^���1<��E�H4 �K$�GZ���x�hD#%�s�@���2�AJ�����ty0��$�|Q:]�F�@���c%Q�ل>�I�4�!'��:�l8�GNh)�
t]y���h�%߄$��V�,L^��3�r�y�3�l�L��3���zG�����������a��|��l����ቪ&�%v��]Z^E}|l|����(.�{��͖_|�ς-������a�\P:��.R=M��q���/���V&R�-�N �����n��fj�IR�D�����.������@�(��M������f�����?�������_�֟zL{$Ꙟ.��7�����oz�;����!���cөd�Rs���2��R=^����v�tc~xC8���H���_�:�ˍ����fvL��?x����P�Qs!{��? Z�y$�j/���$~U� �M�e�pD�����;?�z���]�������	 �#���6D�#��H� 8>)%��;(0��nh?�Fs��\���@���ߔ�~�A����e%��g��<����hA�O��������ݠl�s�r�r)�a�lD��b��ve�qY:�,@����Jo������£��>��>��,F���O�\cՋm&�IdF�iL��� \*�FM��DE���<�����>���+Ҥ��QQ��J�GŮ��i���W��o���~�U�~�����岗�占��4;�*0Ξ/�����;�<|�d4>bFS�zk&�sB�1�/�����T�h�0��r���2���k����y0���ڽ���od�t*�
	#r|���C�։�g��o���?��\��Fq#?�뜃���4x$@���q9%���^-�����4�m��O���[_�"+��aŚF�����J�} ��{�#��� PL�^�;0�JtC#H;P=^C��͌ǘ�k���ZĚ8}��
p`�*X��Q�����)��
 �1ϱ�9,��|��S�@��f%[ۑ�`�S�Y;��E�I@�{Є�M� y�I��"-�]BZ����Щ���8���=
�PqEx�<D��l.e���N�YYD^`%�/�����E�.t+�=<|/�Mf�pIE�KU�4���u`�lEc��y���!��+��n�Ü�d�U�2��T�4����zܦ�I.�H�]t���z����RzK T,��{������|��C�˥|~�կz%�@++2te��t.�Y�{�o�߿��O޾���7��O����"��%�|P:j�x\�zDq.c]��f��3Q������動)�%��_��o�=YȃSn˙�upyyYm>�TʱJ���ܢ�MF��t��͖��P�JK64R�x�����o߾bq5	\���Ď���w���o�{^h.�tB�x^"�d��k�y�E��R�,e�P_��ƟnDUV2�w�(�@(��m9���'P��$0�BA���H"/>�By�$���ʫ�|#� ���z���t�8`�RR%��P'�a~@�	7W�&������^.�jG&\Q��V�kc7*|�8�� �����گȝ���*ԉK�Z>���٧C,�<\#���:D�`X��5�)�<G}�Q�*j�V5K���,�D�G�@��$q�Z4Ȥsl��\����ذwp���vJOb]!ʳ����C�~�oP=�t���A$`���i���vt���/����w���B�)!(��P{͠�`n�?�P43���F�`"
/3��ҥu]���Ou-�wc\nh).	劄��t^$H�F���qF�ie�9ñk��-ҹQ�\���!�pE� @�ʨ���b�L<�e���FV��qc��Js1'368��A�gee���HÁ�ٱ|l�����8|
�q�2���#Vj.��ԛ`^6T.jT�3�S!��:O���=�e<k��V��<N������d$�`���oPHL$`|i�aT��i�P�7� �����m*��ix���o�Ԥ�	b"{��b��]��ײ�mX�H�s$����A/�μQ�&���<��i��er�����AKV�x4`E=�<��K�U�1�q)Ky�5�Y�`Ϯ��Sa�"4mKŕ\4CeU��q&1jV��5�z
] ���
	�&ցTSu��'f�f��Z^^��
�e
̦�Ґj= ���I�(�S�Y�O��- :.�I��C],���Ǔ�z�}v�je5_\�?f	�BF$�*L6�����A�'F6�E���H�_�Z�!����Q:n�'+N�o�e�ߥ��c��T��R�.5rY�	�	m)|�P;��
�IdG�c�)�e��%������N��m�ľ��f⹄��[k^�D�0|� 1�x���J�@2d���R(�b����t*���Й�� ��'�VHW8�H�*u$��C�Fԃ�8h�gQ�(� �L�k6f�Vc�|:f6^Z�Y��-�Z�uiv��]*�GV�-_��Js�sg�=�A��������W�r*�-�g��Y��cq����)�(�&��G>\Ă��d�"k���"��'�|p����`����QU*t*]�Hvr6�Y��C5h72d
��l� v��7��g���?��>�J)�H���Ru���H&18C����爁�U,�p�������v��n�����r�Ѧ���&�X��_K�7V}f-�Ҝ�Ati��^̕�C�2�3|�{�⁂m;K0:� ݾD49��&�2ɧ�	���z#Q�b�'g{k���M��ئ�Q�2�����7��Q����s

���޻��������C�,>&͙�8d_�ZKg�-f;5׵�����q���rP�c�Ċ�ݔ�1����	�����:�C��"q)8j6�b�T��mgң� ��$xX�#y�D"^B�@-����	Յ��S@���U�$�T�K��V���X�.�_����Y����\�	`A���1/p,T��=dY*>����˲�C$B2c%������xnC���s�u��>+k�`�0_F�t�q�Y�%c�Eg�$���I>�f�PpVk��H��*&Ƭ8C��FF-�x�Ċ�dJ�Q�."��Fx���DEc|f����?���?��0$���d��**O}��hO7ċ�]�u�bО�"��wi�N&�����|���������"L�����ܝ���Q��{om5����3�����հ����Dv����	�����it�`��M�'�`�����1�;-�����fa��t�@�uC8{����$�M�D-2���_*`#IA���c�U���R����uj}�`�*b�IGFc&I2l�P"Pl���A(<�T�\e�0���b���B�*ῇ8(22�����v��������"?�)���j)a��+�m9iح��<�P"GEDE�FC��-[� B� |!�����>�J�R-5)*��8��\�Y��$`��x�����9W��91�+�F<�"�(�[��\9ضDQl����K_�b�_�g�2�W-��#������Z ���Nː�<�fX;C�^�k{�LL��!kO�m� E�	O%�&}@����o8���)����=��|j�U�ך�痗��Zu`yxPz��R�F��)��fc�~�-cc
���}����_�����ܹ#b��� Ȓ��@�s������p�%M����y�s���7^w��JE<[G�I���̙�(�Lc�b-��V��]J|-��r�G����oN���<�
FP��%T"�DzS,�����b��:��t��2ng1�k2����8�T�`rf=vnA*c/p
C�t��c|�ʪG�]�?�^ S��.{#�N�f-��6!Qd��a��t�BvJ5�D�VZ�'�1�:,��F�A�X���|�Ʋ�������:t��ա8Mv�N�"˜� L���MѠ�ny�u�Pj�n�j�f���H#�(VVµ��8x)#��qۆ�邉�xC�������Y���8[o�9�	��-��P�R�г�B�D}T��X��j��IJhs\�!�e���B�o7�����7c3r��3�B�_�;KK�z����o��G��|	/72������=���Ţ�̎R���(�uU��	{Щ6�Z+�6��|��{��W�n:5�f҄_������?�;vJgi��SV��eY��3�� L��][-�!�����ɷ�qz��^�Vu2�]JN~�w������J���1ڢy�6J<j5D.8E�	�.�ܔNe��ji|lW>ϲ����ٳſ��O�ȏ��0�:[;����3]Q�%I���r��(�.&����2�A,/�c6�����O9�������č�_��#�Y��� \�z�����Y	���׋W,M)�|���Dtg�i!��ר���`�`��t�\ƈ|�V=]I/k��B�+.��)ဠ+8��a�a�C�X��wgߥ�6�$��L��Q�_q��zL�N
#���W��N_ɝ{�-�l�c�d��:jw�=?|'�[1��z�P�����-�_��R�Q�9������A����:��b����9��t
$�J�%x}��=��-���@T���l�#e�n�j���JE�cW��ރ�u�..5���3E�.x�%�-D.�J�����-������=ik@��5��h���V5N��fܟ�؈T    IDAT�aJ 9�PY�t "@ݿ�v���~�N�m��Pk��P��Y��x5���Գ��l��S�cfd��^��[�u��׿q̊����xH��9J�8|}�t�(�Y&/aB�탻��Ν;�D��\>�Œ���ȁ�ҙ���*S"t)�p�d��I��"Y�
�Z���;.��� ��F�vuY<Z������� K��'e��s���y�0�YȮ`���ϋ�ٙJ�gϟA�`jr'����>"���:���Ba(��X���y;�����x��%��:���8 ��2�:#�s���V�|�)��((0��mп���m�Ű�/��k�&rT���JCl@�z��.�l.���Z����RM$A�%��G���_(r�b�B��ݧ'��;���W�>�����{54ۡi��2�¾�k�q����!�K�u*v��Ë"��	�ڐa׬��hi�۰�QR�,"�v!���I�)#�f�����9$H�OD�φQ�}_,l7VR:�z��F&�Pl(mFA4��  ��x�>�Ж+�4"����8�HLyJx-��>!IЂ`�R�hF�[�Yltj��je�kű{G�\�^+��V�[���pš� �e�	
#�T�oԗip��h|cuuE} �քU��%�o��&�5&n��B�A�B˦3c�b??0<�$GP|B=ү9j�eeBY�\�+:(ɤ���(܃�a��~vtW6?���*��F:U�XL��D�����W}�w����PL�)��I����� :����U��˴.��l�|�m
#HtsU����b��J���'�Q��/�^_RRy����?����]�G���ݺ��P|)i�G5'��P�^ҫd����6;l���@'ȳ�˘�G�5G�~��%���:{��k7�q�L"��y�u��s-�ϑ��EV��Y�����H�5������3-��ݖ��W_R�z	�%���}E1OQN��k��y���u�Π7��Q(HC�PC�.U+�Z��v�͈[��Os)�H%��'A,�X���y�e�0t���ܞ��^<^,-�q��eS�R�R\M%Ŋn[2�G�M��<Α��<؝�,$?�C��x

�(�W`F��z�_:a�p�Jcթ:݆��<���g2�-kF����+R��p޴�+�믹��/x�W�b,a<@>,�͠k7U�t�p��W�����P�8nY<{�������]Z*2��2A���TZ��m-��<���^|��u��8`��_����|	� N�(#C8˗''iV���BUaî��
��|�o󑯧:����QO��,Z��t���2�X����V�L_�t5�:-���wTh�?�EY׈,Fa�-p���HV����L)���o�����f��_ݱ�=5Q��l�g���Y��1gj�J�!�!���V�����IA7�꣯2��rYD���ݗ���Q|<�LM�Z7�-�F��0Ƥ_�߶�֨�M^��{�W�hR�=�E���� t�<�/�;��,E�x���B���c�p�װ1sb���['ru1 3�|
��h<� I_^-=��Cш�ǏG��q��E����)+gFj���e�$Y`A�z��P�WG0��2l�q���-/��J����4>=62z����Uh��tŸ ���\$U_ݶ�'܄͊�)xB�jb(�g�}J�-��_�����?��O�Mk-��t�������zKШ-#��'<�S#�d�Idaٻ��>����<en$�ŬH:���D�w��BK���Z�C��EV9b���3q�_6�bzk��2;�0���	���L'���-�l<jbs��%F��jD(��rBCo���
� ְ;�����J�2p�Z�Ϣ3��E����2�	o����%�J�uM}�q�X�g�v͉�������:�wW6�K%F�e!eZM��!+|E;�<+k0�œ���ODC͉���L���?� zA���;�%H$�R"0��T��1�l�5P��W�n�~7�~�|Eq����"q.�2ƥ3#(-,���wd2�����z���G'#y��*I��S��N|;�x.r3e���8�Tp���Ӌ�Gq�1;��%1�����#gu?fAԃ�b4�M�BNED�v8mU�� z�СCG���iqanqqaǞ���·Zfl��
�4.��O#����\��I_���y��Eဣ����! :�{Lf�j�\^e�(�	U{���ࠚ'�#"���X�l��~���ТE�7a�b�
.�ج�	������c�Z+瘇:am֔jwc7��j���;ks�]������/�1
�!+k��ե9�LO-Vti�X/��n-��ƭ��o-��x6�冕�A��t�qX<��!��!���[�3՜㲳���a6���ٽk��3g��]=Mvf5j:�R�?̿	.���n���Պ��s~2���z��n-0S*���i���Q���ʱ�G�L�ɨ��.i	�-��ͷ�}�-��É�����[.��'����Ę��<�|؇ߔ�""BS	8��d��j"��&�q_�4�tG`;Iaߊ�4�]V�L�}�b��a�D[Z��9ɀ1���D� Lr@�ŒЊZA����{ф��E�H�F� ��M�z�dC��dEL$%�(� +�b�C�i�coQ����h�H� ��
[��Y�E\� ���;�6�Б(D8��:l;�?&f$FbьkN�M����PS�e�oc+���ͺfm�u�g�eX����F��s���`�&�e�9��C�Q���tX#�c�a*��)����F��t�)QZ�T��`X�� C�:����^-�U(	)��"E��w�\Ħrk+��N�t�zGڶwN�����̣z���%l:Ryv�Q֗�⃭�e&{q!5Ĩ!�NO�=p���~����vO.����Kh�f��:몃{�s�M`e�=r�/��� !�=X�@�d�-�����E+�L��Hܱ=��V��P���=r�Ql��m?u�Kn����1X �fs@G$��_����hX��J��v�\t ��(�(a��7X�������#X2�A+\�7}L31�^��)w>�@ּ,�r��g��^Bs�-j���I.���Y�x�4Z��B>X��Y���}��6a���|�!�k �/d�j�J>7�b��3f�Yff��p�K�>X	K���d�շ
��O�%�#a�k%d��F�	[ v۲�i�(r��,���K�d��+�3���1�Pv��x�Zx�R	�\+2XgTl�4.;e�� 䜊�Hg$s"i��4��i�+��j
���K_��?��[��j?&!��j��1��"�r�L�x��E�&�
�``��Ot��By|�Gc`<��oþ�����g�G�+̚�wX+�Q��&@X8M�k_�����=w?0=݃K�L�tQ��^�9����##D��pZ!�P����k��;�����?�Wx�݈��w���eK�@n���b�^�Դi��,R0jB�n��!�}��o��3n��֗������ӓg�"ڨ����&�N-���3e�*�ݙ>�6�\D{O�8�lD�~z�������3�3���r��ڹ�+�?=5)SoT�-{�0����=��Y�S�Ѭ-���P����"
2I��a�ԯ�z~��\o���H�ٲJ��y��i	K7�Ȣ	9�h��d�1+��M?�h��7�\a�-VW�c����.ߛm����a�c� ^�L�>J"��A�aW$�H#5�;.̝n������S\h��|��1ۮ"�v���y�� \����G;`�c��-���q�N�bc�;����-lp񝇡3�0pTW���Ȅ�E�U~ !�D��^tV��a`�梬�?��8�p��{�\��gްs[�f�֘�ʺ'��I�W/���\���ݣ��.�wWx�})�m���߅�Q�/�˲�̜����E�jĳ���ml�'�zH9{m��N�����5�v���r����Ęn5i#����
ĔT��pa����x��e�g��I�RA�����ǽE
����s'�4OY���6�f�^:{��c�3ӵ��˧��T�]j��<��0�dh	٥�sb� a�􈻡�{�o�[�P =qpQ�d��r_+�a֎dsW^sm.��2����ٜ��Լ�^�0t,#j{%�*�J���-G܇q66��8�!�g��+�8���J�N�L6��=��w�U�Á��`�όF��,"7E]!�������\�sB4��_�S;�8���=/rmܦH�B�PF?4�^��.z�M:�eV4ia>�"��)X�s���Cٶ���t�4���]��@�o�C��dD�K��7I;�{��!�.��b�]�R���7
��6<��H4��A�RzD7H�|i��t�r�*nJ�*�+�d�ݚI'vLό��2�z�ٹ����}�}G߅���]�3	w%�w����qth�C��g�a�Ӥ2=��%�����Hu݁w���u�s-O�$�v�=k�����6[oe8{�X��3m�hjF8s1�����1����e��qm_=6I�!�'��X��9`��f��#���2�a�h^t��+�1��O�4�b�$<z��t�#���]�&�r�Đ��pP�#��C�I�9��^���6=�Δ�U�a�T,1��H�v���hS��6�C�
�B&�R&�|���^�����l��_G<F��K+���*<w��m��A]dd**EKH�K$�N	���5M�ً�$�{5V�W6"��`���"��#�W"�\jff�t<j�R��CA*�ʺ?:2��mQ�1PxФV���峆"�ZR]�L4�Q�ܱ��sԤ���LN���)��y�� �(���Q�t�dh�ӏyk+
��ۙD~����Je�:Mf���d2q+��g@���:Ω��=���
"P#�������h�Sf�����G���6��"�?7����ȶ� <�&3�@�=ۆ��=��g"�gˤVҊA����<i(t/C9`bxI�+���������'�A�b%w��'e��X6E�l�M��q�];r�.�ѵ�"W�ED�#�1'�":���E����؏J����'��P�x�r]��c��|�A5i:	��Mf�\&�T0i%0���4M'_��\���5���;��o.�xA��r����i8�zU6�Ff	��T�2%�<�y)��#�qѲ`�Jh��잙9�h �������AK��p]�3�a;�!�=�p�gK�*a�	�J���^�uV�8�qg�s����+X�$-L�Ë��?|⁇N,1���,�-W�$����e�;����T��_ ��}�n�og�AE-��T]�J�i隖�_�5�r��GІ�{X(��%Yq��B�/h��)]�A�Ƨ��0E�����
��L,�vha�
Y�&9��FFr�'[��Z,��b��t�
X�H�� ����/Pg(��DpQF�N<4�rz|��STd,`�@镐x��Ag�L���3ܧ�/&9���H���������L˫%�V(@�ӈ��1f7e�a��*&�����W���,V3�N ��Nc"�@s����(z��!�0�t����1��J���W�T]Rr,FVvA"ZZ8q�t"qd¹�k/�b�tш���'N�=s���s8��%-��-ǩ�Q�� \�M���2��Rڵ�Kr6.�|�B7:D�a�Bz]2���ݔj�Z�pW:X��L�O�K��s�~�ޕ�!V������K�x33��m���}����W�փ��֙�ŢY��h^<��Xd���F2vde�A�zX��T]������KQ�71�iX� ���3�|!m$̖_M���Hxy��s:�y��_���J'��2z���s��;>�w�>�|����Jqb��0�SG�)b��*@*.����#�V�]�[��qΜ��Ue�R�nʘcm	�+�b@+��ƞ����]E�GvO���J�B+��)������@�̋���EjK�����a*��k�݀��p6�?0��� `-ڙ(uB체	��n�X+�@�[��px�2�I�CX䗱�*�m|+���H�:m�	� %�r"\�D��@�ؼ�Wa�����h�֠$񄕃%�T��e�6+�&"-� �	�[��a�lˉ�S�o�B�4�G;MyD ?6��_���I���#�?H�tk�nt/��H���Ȯ�[�y����Y�����[�u�5�\��J%�`��<����*�G�<F˷�Y&�d275�{�Ƞ*�
3$�,����t�K�,��_*�Y�|Tv6�9��.@�(G�4���܎�*�
�@'��!���{ <��(D��)����n�:)��3!$~�)^4:���"����L�2H�����\blvA���T�0�bke���J�dZ X�7�:�\���[cC䥀KAb�? (�υ8NA�������t:i?����S?���?#�O�����¹�g��Sn��9Ͻy���x�K_�k��{N�+-gQmA-qk��
�B����*.Jm�����OX7�Y�?���&�Z>a�L���=R��`��:�+�a}ZZ]q[�u"f�q+�p1�k'R�R��0�@�v����
U­�*�򽆽R\Y�L�mۜ�]`M�)$����yИv�{T:�ǃ6��Qo�vs�$��AQ=�+{�	�=s&�ȡ�+���i<*��=��*f"d��d6Q
�8����숹y��i(�|�i���ONӿCM�l��]�Hnd,�H�Ė��*m/��k
�5����!@�	�L�(K�\�&��D�	��0� .5����?�a�{�`
Y;8\n,�*�p,�-&�,&������;q���S&�g���_�bc'[��J�2���L��Lalda~ieuI��XQ�v���zKM��GY��O�o;�7�z�;:�ų*�py�����E�ҵZ6IfN�|k RS��S��ѤG\L�տAp�|�������|Ϟ܍7�899�ģ��#�b7��FB��,�^�eD�P���W,����z)p��T���jBxkdֆ��_�o�JKf|��I�Hqد��f�6����x˛^�co~�Z<y�W9���p��1:e����g���������_�[8��B� ;�G�B(.ڛ�E�Ht[�x�ź@z���t'��f��6r�-�*�$1I�$���8;��`�o�����������O�R]J~������Yt��D��+f�P��#�ǚ*��Qm�����W���dg�kNu�x�Ro���v\6Y-�8��J�B��D���)��f�V*J'�-���߸�v+6)���j����=z���{'dk�Vy��[זY���u����#�<#���F�Z?����r�䣷���Ǐ�񳳳v��5�tʣu�2)j�Dq�wp�"��H>a/@���}ey���-y,�=;���	ї���f��0L2�XCeU�E���`&��痊+'[^1k�oz��ㅝǎ~�K_�z���õW^;�ߑ��w�طk�3���-���F���?8�c'���塥��\�Z6,7�0߆�U�\w,�koP<H���,+��� GNX)�5�9�48�F���Y��@�F0N�����dCG�?2˪L���av���;f�\}�S��D���I�,D�NB���i+��؍����OO�^	U����Eݗ�a�IJU@���/{�<������}��nR
`�EQ��X��_�^�s���W��_�z��#���H�n�RO��i/���k��������\���S7�㿼��l����k��9���0���
(X�:�P���G�Y�W�KtO���S�!�e��p����Tt�9c����{ �u����:��ȁ$���LQ��if��<���c�g�ښ���r�k�ٙ��vg<;�v��%{5��,Q�ER�b @�����u��9�������]���8l^�w�'��?���f��cG�G?��̒H\�'�����Ke�=���VW8�;��re�@x ��R���߷d.���O=�̯����R2��p˾��½�9r����݈Hʒ��Y1=�EՐ��Φ����SO=�7�'��>m�    IDATs���]ݑ�9b]�~�D��R*�!I�Q�~.�
��Ji�*�+�`rr�СC�Ģ}�ji�ԫ2�-$_y��cG�����P)������l5"QT4<����
M����5���1���+���_n�<��XRn��������U�]j��������j�+�R�db^����Y^ZJ�r��R:�*�	�@�	r(�G�n���B"��/
�	Q��%
�e��4cD�U��f�E�ڜ�M��峞T���aN8�	�A�7`o��-}��`F��E>�yU���E)�u85�9I�1j��ĩ��^��@{���0�Jh��o(�Ju����zb�@L�1�أ�$?��P�e�������!�JX?��ݣ5�P�!^rjvf4Y�TSaOӱ�\�#��>��?�������3G&�����C��;2X)@g�
���>�ē������?�D����7����?Ǵ�2l�t&H<��|\D@p����T�¦Pm�� \�;��:���R���ٸ�`�XW	����������-�݅����L<~��xR �=;�n��`�
I��<d�͢)[uT�.�� 4�;Jǁ���\"G]�,�HX�z)���d�eۮc.eq���������s� @�*IN��=C���k�Za1�4_K��Pl���LA�Y�JZ�I���l=���ł�ه}uqg� ���0#�gU�=��~p:ZB�׹��>�Q�D�����=ǉ���d�>"�OA�ß�b��.�Q�p���m�����%���Kc~w��n8�4�;}�AV+eL�|�,���h[V�يB��`�K�*BK\���2������p�.� R��آ��b=��xw�X���Y_*#�H�D�@�H�S#Us뇀��P��r�Bm�38�W��[,�T��`F��8@��Lɳ�[	��"_鲎�`4VrU�!���������$��ځ�&`_�a�k:����%��d�|*a��X�uؠ���rE�a���	�G�V��@�l ���E����lj����][9<-�΢(�e󾑭;<>�CEUq�r�o�[1ffC�+������%��R6�p�,DUV����F:��e2�X�P����@*yph(������p�J����?u6��B�J ���!�8O�5*5�Y!E�J�"r�b�J�i�8Ml-��p�^&�6'A뺩�zm@���P�P( ܆jߦ�ؗ�� mK��􍲅q��}����T/����v�`�	W�^M�f�+ Zނ�k(n��A?���y�e��=��ø�C�	��� `����c��Lg0v��`L3��j�RR�ʀ1�>d`YIB�oB��~��>��i�&ؑtt�� 9�g�Ll 
ہbƓ�F�F6�b��S�xqm�C_��ؘG� ӆ���tY� }$N�g����?��jf#���0iB���u��eƟ��s�"�Y��|8��f�.�W�U浟_:e�%*w�{ V������]�l-ǧ�K�@0v`���wT�~�\>a��J���D\�K'O=�.�>�o��������=����F@,�_�o�~ˠ��б�%U�f�nx!���f�J�p�=
$���"�Ҫ�z�%��꡵#R��o5�J:(	o�/�it	�!�A�r� �����[��^�����\�����?�4 �E*A/F�~��8�E��6������{1���M��!}�pJ�]���G_�3�"~oe5��#�����8�a�0��?;9;g��q�G;!�aeBZ�d�J��C�:��Jd;J1�����������c~f�!���X,�}���2/t�-�'���� P�Z�`w	�5�A#MO⚗�\��2j�`�0 �L�
�ȉ��&���k�A9��<udm��L�V�-u�F��"<�ޖB�dc���2�t��@���ʨ<U���H����:���>f���2r��ȭF�?�XWP��]�`϶}�ۏ�&�H����m��h�l����������O:5��$�(�PS���`��j�S�[4�#N6����q">�  �\IDO�	=����·f!�.!q��,�?����t/���x�"�y�Ғ2)A8�\A���_��Ͽ��y�.έv!5�#�U���p]!M��j���DN���`$���8�ˉ�C��ka�ػ���t"��څUs�Ϸ�,q7=~l���^*e��i��Qw$S�����)�ɩ��Bhp���(�5�ff������w"3���r"��׾���9r��5�y��H��*�%�8!�C�F\];�f���M3��l#SP-��@Ao̢Ҁ~�ӹs�N4q�����$��Y����������Du"��.��m۶)^��:�y��j�(� ��o6�m=;�.aF���0"�/R������q�k}`V�i�Jky�P� �w�B~|� f=%W����qYKLϥ�r�ص��+��v2m.܄#�-���� �j�xt��DghtS C�E�h@!�K։���DƽU�-V0.U�R�NO�铟 �ƿ�(��ҥ��!�aGI|�M�;�hx�V�}�~���~��ڵs���y��`W@��)�.�|ʡd�<��d'!"HSA
�����.�]'Gu��r0��� X�����v���Fi���1w�q�Wf5'bz�p \/G�&d��&pv�l�/�V�#�0�NBf%���`xd�����ٙ�	�'�x��ӭ��H2���Iwt:�8���d�V�D��U=}���O�C�����0F�b�9����z�!�K�*�@���[����5ș��L��t ���S���[�Y�vؙx��fo��`���	Ni�ơ�AV4gm?�yt	[J	�Ȑ��) �#��5�.��&Ϗ%r�]���T-	n�X.H�#O=����L����H�wԹa�!��
m��1X,���22�Opͯ[ť��,Q�N�rY+�k��U���ID�`���KOW� L2�<��H��A�PO�Mx�*�"�"��6�9�#XN�TW ���z��r��Ȁ�j.?l��D|�ԱS����@���WfY��;E��_W���JP���*T�~�݂=5��я�HGf�&zG�)E.�c�g ��wy�0=���(���'�QEt.�ms(�BǪ#�O_dA�7	�?aRj�h7�G�O�"���]��>�����FpGr>�XJ/��;N��>�ϟ?ϓE��%�UW�!�7�4��ȥߚٮXD�@F�L�bH?�add��������!�T����:.C�?�W'�$��ԯH�9�S5��`�A֌0yh���sm�[�q�.ծ3����O�<����-f��	��<)b����<y.�\��F�8���'N<6�)����W�
�,!]8~���cOF�Eo���M,�g�0J�;�v7&���%k0$n���Y�B620gr��:�5J|e��%��47F��������!�H���@�t��+�-��Gj���P�6��!��H�5�ԭ�A��z��J�9�8A#2/΅8Y�1����]��z6Ł[�>h_#��YA����������$2S�d��P��!�-J3x�_�6�z���2`i��/�Y��
�K������_Z�t�#������v{��EX@���A���@e��8N<�劳��kǎ�[v�M+���X1��	v}���Y$��繑 �CAy�(cu=���{V��>�.��sώ;��8]�#�`S�+BW��4��O��:B
_�ͷf
E1��F~]q�ym�+F��j�+<+�o5t]
/R��K
0'f��NO�X����\~t�ޞ������_�i��֭�[62��b�i/���/ν��޹��{?07[���{��G0������YEC���{��QGA=m s��	Ę��[1<5��h��n2)2�����A�DHv	n���X��Y�%B��C��Dv,����*�2帪�<i�IO���d#�����$�{�̾��922Z�r��}d�8�E~�"�H�}�zQ��=Ȩ"lFa�Z־���rJF��47p�'tj�㉱338�������L^G�S�D��������΅9�\����������#c�q�^2R�����;����l�)\�A�����
��ؙ� �Y̤P?U�-t�E�%?i��enV��g���t���j �f��}�o�@B�W���X]���L��х�Ot6�4u�M]��["��J:qC6]`�ѐ2��+��e+~�a����a���-�1�t�=�b�p�0�p�K9��6�A��I&���������;|��m��W�Z���}o$<v�й�W�����-;��������ɩY�Y�0w�XsBX�ꖍK:cG���|��hHt��r��qk,�[�U\ZE!<	���%��#��d�WL���tªzɩ�q!I�Pg�	�Ҥ"5�?�,y�n�)���a��i֢��'�� ����!����Q GG���/\�#��(����Sh(uE��]��G���_�]���T9BoN7P���B��_=���oЮЛ5���F�2-&p�b�3��c4����~�?|�ۏB]@@4�E�A�O6tiP�VE�h�Ju��[�͒�A�7��]�/QO��,������ٳ˽!Z$A�[�2� J~���B"�h1�	(�K	�Tڬ�?���f5/��W�aBuk`���x�#��گ"��+����Ѡ�Z�C���|�B:):η�Y�=�+CD��R`����[����)AfB	��r�t�|H �J!'A�6��pG-$�O��֝.�){#�~t��,���-��⏳��|RTo��'�����g;v��y��ݷ�7[B�L88�c{$��1�pl��??����C��v?vи��h�s�?�ߛ�j��WI��<��)�����������}��[4��3�H5�"��t5�̡���R�`�.��O��q64�؆ȥ��!��R)P>8���~���f�C :X]h�LD!O��BوF�08�q�Hf�eun~�Na ���o�;1>>y~r*��bySKT/?���y�1Y���aµA���!T{9��C��\7�wt�閽_LB*�� Mƍ�0�F�lp9�W<B������)�)��P�R"��"B]zhؓ��O���W�-����U���Uvvo@�G9��,=���R��864�����C�o߿e��s���K�=;��{ێ���^���z�?��'{r�RpA�:���/��;�.�����}ԥ��`�2�����39gN����w���	3׿��I,�oݱ��!��2�Ů�CT=��K/)Ap���������V�!B؍M������z��Cf"l��=�ra��I�� XP&��I�	+ec��ғ'W�xL��*�T-�6+u�|6����P�ӟ�@8���c�����X���$����Lg��w�%t�O��@�^�|"�p=��"z��$��$O}�����ܾ};��8���Ȉ)0qNX��$?��!�9<�Ꝇ���d�:�F��%f�+�<���L����=қ
+Xv�6����<�87����ܽ�lǐ��[��<�T=�⡗�����ȏ����H��\HN`3WN��-���з,��j��щW��v�Ū��h(;���ɭIq`�VLA���Ǐ��ٟ��_=���=�o�9��9H�������,<��� �E"�f <��檤�AL������ݽ=�4,.�/'g"Q��>��?��-#=�b�R�"d���ؐB��l܊r�W���j�A����H�ܐ~B�B')�Y��Eo_�B]ݡ`���Oq��1J�p�^�ĩT�B��:�RF�D���ּ�v��Z����#  lE��@7I��e�NL��Ux��I���_3>|�P0Vd 4�l�WWB��@if�'NfHT���ϰ�� ޼�C�yt�;P
+OhK���S䑫%�Ϗ�깩��qt��\w����0���Scc�#��N�<?7�)W=�����3��D-{qAؚ/w���ڭQ����*��4PgWuX<�@]�	6��C5�������S���Ы��ՒG�=s�8���w�aV���@��(�㲉
�p����_��f�{����x��Ƹ�΢�SIa}����F6o�2�!lt��=;qא��X�B|��Ti<����F��9��=���)�(̨
sU����d|~~qa��\�$�
g��~"TA�Y����T+�8)�ނ�>�'a�U���W�t�Gݠw�	�l� ݧ� J,���}����'hL(�� �C5�d���Lʡ԰�NC�q��Z�a''���8v]�ˣb{�)0+6z|}C8+c�0Q�]�>:�1\��s�=�X�WD�"�����A�x\>�pW+y�����c��1vM�j_�}?R��/�%e�I&�V�(��Ysڜ��s��^x/�Z�oSgdX�JrR�<�}� �~��T��D-q,�� ������~;66�]�x���	�0C�	%�g�J|!�bA�;��*����/)D��V!'{9������]�b��,bD��D����`���[vHDX��"!�eV�Fy͈�Ćju˃:�3�� 6�	��aW��&Ew=p%?Qjںu+�mbb⩧�:�<h�̙3SSSd 3#F��f�'e7M9��"���M��w�/6(XX7ͼ�3z�"�G�NQ�A@�fl�� gs$>��`�Ή�lG��V��ٓ�X�rG����W�N𒚷׼5Ln�¶zeI,:wjh� �	�Tm�c��B�V;��v���5 Z8�r͂[G�L���ž��Mw��B���8���0���d|���?�����a�/��x:�>�K�Ǣ�σ�7�W5�t��x ؃�ۯ�:���o����b	�5�X���g����J	��J6���:�$"���F�`L"̩~4��Xt}�*�J�'*�I���e�"��X��sc�/�v9B��Y�zgFH�'qf�$2)z%����eO~�X��u�N��h�HD݄����k\v�+����i�N���ڌ2z�x�<|B:�D�]O~�޽yO�0�|��ɕ�w]*0�� �*�6�6�f�Y<�[�$�U��U�N����Q��0��u���kB�ßJ����@Ѕ��	l ��l�qM{�qG N"� [�����d,ڇ@mۻ��[�8y|&���n�{�3�S�P�\�ypF"v0�r��j�V��#�%*���[�p���] ��#zC�@8�_ʥS;v�ڌarܜ��L�$St�%��bV6ą�8 l��.`	~%Ǝ4L�ő��$.(��3	��܊(�se�j��W2)TiR@j�h G���H'�O.n�u���Anٲ�%8�-��'\�[�(�',�g�y�����9#(;�:�F	�k��j���'H��|J&&8�Қ˿b�Σ�Jۅ^�+��y��w#�Zw�q߼4�s=~zbށ.Pئ|۫Ƣ;�D����6u�墭��+��/'�+0h䱹�tY���(�Xj�c��ʈ�#���oQY	�������"��}��*����*���Xr@ ��2�3U�B��a�6g3��̟f�
���j�5e�P� h�hb5�.�9-�3E�Ϻͅ*�Z"*ʩ����.$J._yva��;�t�����u�]�Ν��靋��P2o�����3Ao��;;3�j13�`&uc6�	������Ԝ����c��	��9�[P7r�{��/~��
a����,�r�E%�_�Ƞ�J�S�֮�V�B ��n~�5Y�p�`�"���8Qz/�#G�r8zD��Rr���ӗ!
w�ɭ�r8����Je|?���q4�P�n���m�Z�8�/#m[��ɸ�"�^Þ��] ^������:⃃���9hC���8�SHҏ�����FŞ=��� S
�d� ��@�B
_�(���l-{B9�m�۷��`<cˑ�Ju��~R��qMo82Lm�ETm�����    IDAT�� �K%��2 ���I�z >@���R���b�O��"�'�0�ZgQKL(����p�&���:䞩�*j�Y�d�nw�k���r���,��'��2F~8�K3�a����Ŏ�/�,K)��&?���C*NV��|%��Z�m�T��?���A�Ja�(G����r�t�v$���0�-/e6w�=������J����b�ܞ�,���vC��k�x���/����%�kxs���w��x|=�1qe�9�;A�9l��D��$1Y��@0lZ�l�o=�Z���G�:޺l���:��K>Ag�;� �����h�a�ϣe'�F:�Kp%�E<U<��#/����P��m۶��[��ƛd���|�b5>|�\I��d�Uf�Q�"w�O���	jB���A�͐mӖ��N�׸��-86�_w$��%&&���./�/�(��Z�£wa4#�Q� .��g&�0#8�qr�e3�0G0����*u���P%Q�i�;ߑv^�B�f�i�$U��e�.~��fO\֓�W��Rf�j-�r����L&�H����o(�[�K9�@��Z4)�ҡ�s��{�?�Z�n��w'�YWȇ:�O:��6�z��O�A�c`�'Cd��a�WK.���W����hv���Y[p��%7�ou@I�&��f�O��:�G�p��9��0��z� P������a�c�֭ �I{����l��y��$��ʌ�C:��˓�f��<�hfnO��eQ
���!�S�g��J9�d�a�.ʯ)š2�Bah$+8���R��J��rLjD�+�`w/���,�!<�"|��!0�q�jC
4UObd��{|�S�鮖�E�.�{a����z�k�X�b�t�'u������E9*���L-�*S+wz1����w�|o�o�rn2*#C[ȃ|�2Ć�n� ^���>��͋o�<�(x4���rR�Aε�<��Y|�������^t�9�� 6��x�uy3tr^�I�(��@R_|�N5\s���V�i�-y A���5)�� Jnf�6­�(�
2'�&�`F(�
��)����<��W4��~�nobΊE�P�<HGD(��� �� (C��*�jQl���q#��K���t)�z�I�O%�!k>�'��s_�|��\bZ$�#��_�����+�N��ӻ-��������7�D���6����Z6�
\����O���M�DJ3h^�M���iֿDAh��d���$(�x��%q.�JbMj"��#Y*&��L%[D9'��'�q��\��ʥ�'\�s�dGO��b�]��B��0��;_Q��=#r�ȣW�X'<�-���u���x����\-C��X��ռ[����i*4�N��AXԪ&H��}�z��$��<|B� J4�0;������d�́O)MC>�z(̧��[��2"]8
�@ݼ���� H�V��:I+ ��P�\0����+��v��n��hO��2"3E	w�;O]bCP�]�l��DL�T/\s���jey�|.==2��w#�D�u@��?��G��{�� ]���R|��YF�E�m40��t��̺��e_:EM��-��\��Y[}�Rw7|i�y�8y�PJ�mc���W�`.��׊F9�������H��Y��I.��af�s'���=zt���l�������'��B�eՌ�-�cc���N�gg8��rzs�[kL���ͷ�# Z���k���˴Z��=5�D��$NY�|·������1��4����d��&@���l�Q�K��R ��L�ز"�:�dʾ.XH!"�1@��@%�\��f����'s�Z8{����=�
tS���R�#eCus��YI��ܮ:������s��ҙ�������s`ۮzz)U�zФB9�-��g��_���ͧm���^�z�S��}�4Ɨ�_����Uh7]��B.�Ӫ��C�%>����A�%JA
�a�Α(�yk'O{��'����d��<�&GoW(TN�x���}��N;��'0J^d�Ky��<�_�`鏕sY�[�rvu��e~�87?�̏���^������Z+�1]r���q�)Mx���$��Or�B���8_AW�f�OAv&�kƉ$�v�<S�&0u���O�l�mu����h	BK�O؝`�	�漇�|~���{zpq#�F>Qy�է��.U����l�@�"<����R>�u�>��������3ScO/-�z{6c�yy��;����K���O�W�����w��Ŗ����zxX��:Sgw�	3wѓ�eU��<�)V�?fr<����k��M�J�5ԯw���Ї?8u~���G2��}�� �����c'ǣ�̹r8�H+�%B�}<0�xm��᪟:s~hh Db�D"��󹙹���-#�X
���E�j��w楉5V���<����`4���H�!p"�,����S�����m�~�4����ꫯ�1A��6��I�`RJ�X�.�~Z��*��|Eè�l:Bz˾��\y��vU�c��ԝ�+E���(v��w�zy�lػ{���M�(���L���@]�n���B����kZ�,�*V�pc)$���rΎ��B���;���~�}�޺0wx)~���936	���Gb�@�9�}���gñ��_<r�ԑ� V9����\���I=i�Ch�d��ӛ�k5=o����ʓ���-SM� @�T�a��2�V��D�/=RAJ��v!3��f�z��<1HM	�1X)kDԜ֊.j�{jDH 
�J��e =R;3/���T�`�{��dI �89��6$��o�����Ӝ�Fw�h1�j	�6x��G��%�+�P	@��r��uN�U>�%�4��r<�>rO�8á�r���/����+���PS�*.�tHa�?I!���ԇ�N�qA�K53����T7�Q���H]�EO]�EI�X�H�U����_�M�ٱ�ZE��O�L��\� N��f��$2s�M��`p%?5:��:��͖8��pm�P/�_ב���W��\6���>;}�����r�(�@��~�����*�A?73yn��wn۾yt��;�u��O�L
���qG셻qhZw"����Z�D�������?x����̏��e�v��޽�FG�q���Ο<59��y�{>��ϼW��]r����uH��b��q�Ɵ�0��~���24�k�l��K S��~Va�I�|��?q*K)Ԣ����%E��p$Ն&�8�-�r���
��#/j�rr�z,�O�5���>���������[�m&�} R��Uz��"҂$��5�pֹ��c���`���"�y�߃�\ٍ%�<u&����{��E�4���|0�ڱ���ڪ^�If�*�H����}�*
�R$fG˜����,Fn~X��˃ !�m;���})X�:x���|�c�޲v���j�R��5A��o=����s|]����V17cw�9����������׏������w>�(�b~�������ر�|莧�y�?}t)~`�n���z:y߰%r���F^����M��V�A~��y���ԡS�q���0^ �H��&�;�n'M���/D����,3�p����%��� @�\ ��~_�V��/�{��k_���z�F�g��K᜾�#\~C�
Uv=s��R��.��%P/�3�gF�CT�"�g�J��695���/ֲy��l����R�:�L�a"�ݼ�2����%j�9��*W#pp:`&�(5@�@%��b��UU��*U�+�G�U��C�\<�����?}�-�z;��\ӗҋ��yt���Е�hP\�jd1���߿��߻u�??}jz���=`�7�r�0�$"��B[S��^:�J8�U����;q�����\&[��p5�`=u�����û�!�0gV�	�ZT���V�>�l;<u���>Ӈ�f�*�2_�-.)$?�=���E�a	8Y�\�@��흙�~�ɗN���c�#R~W+.�b���)���H�wP�J�c��S.9�t�aM��A�����D#��D<�K.&�˕Ztx;|-%����Х?��%�|�cd�U`�_�`^N�u�d����������I��T����������''���>�Ζ �j6������'���N8�1v�22@) ���j��H��48=-"�^@yt���۶���ϡ���;�ѡ����ƻDP�N�sہ�p�aK�L��_�;��y��-�N�t���C���`I.�<}�<�P�X�\��[0��'`d~�����Q�(@���p�e*�c��.ET�Q��Px�9]B蕪.��b��V�2
"�B���05YA5���J[O�\a{]�-��`e*�M�<h݊�r6N4��c�	��՝�.eZ� �8mH�
��:��q��QC���}eqքu ����an�.�z�(�8O��v��f~s �1d$��聵��a7?�ʼ��$��tq�I���ǧg�9���b�T����{����j%�Ϗ}���~�ã[�B�\�܇0�]W8G��ΣK��	_����6!`��Y���-̽�����n	��:]�5�@�y����Ȟ]�'ξ�8&���tp�7L{��"�,��^h�\,'��.���(!�@��F�E'��#�uD-{&�0��u�A)r��50#Wg���R��&��.s�j ��v�69�a�l���VCA����g���2�k��.�R�h$��гqS[[A�*�=&<*�aJ���_�ڡ]�R`�!pL�b� �=����TZTh�=�N���ҟ�᭍ #i����iF���W8>��M���*�ӧ&���b<����:!�7�E[)�J̖��Ѱ�_���>��n��1�X�	eC W HW��G�U.�d�HT��ʆK	�
d'���`�v�-r���ky\�r�_���S��e8q�q׺
�j*���ò9��b9���ғk;p��I�����p�A<�0Ӛ��E��MY։"/�dA��
���]B�3��/�]��@'�e:ȋMN�4��C��T*��'��V���7�a���߅pi
N�^�(JNZ)�R	7؜UL������Rd�VW�'��ꡈ7��b3�Vsxw{��R��T:�0xӸ݀�v�hQ�#��7�2#V���cF�2_��b���p:?�>z����{��rT�^��!�R6�T��o�e�{�s��~�ˀ.�y�N����"�V��XU���RcŇb�/�PV���[^N!bi�an\�Bt%נ��s��EY��T<���)�Y[��?P*Yg�����&@r{��kZl�+ٻ��t�?�CВ�z��{+OLd�=(E�����K_Q7��U�!4��!J�	Z��
٫$�`/ָ�]R�ɍ$�]��pd�a�#�L��10<D?��l�b2ݨaA���K�Yc�O�@�B�T�*�p��P�k�#�	z��~��d&��)k`��U`�t�F}��Afg�Ca~kF�e���GG��U�*'6����<ʲNO����>�V
B�E��w���?���E�]t
��,�
��o>B�T��(�z�3Rk�8O)�^���([�[9�N���F��ܹ��[ax[�1����Zj���;vm�	f��z�E?j�����s��n�+�G����>�/փ���c�����w{@$v<p�"�w���jݿ���]�s��k3�����E���PM����Uß*��}��#����FO�,��E"���SPj>�yP��}�o��'��2Bެ+�O
ݽ6X����kE! �K�9 �w�/���xc量<s����(24��w�ٛ���	$JQ�p��}Re>my$`�@gbIO�j$Z��Xsc=��E�Ƣ���E|�^��G���)a�0�͠^ճ���V� Ea_ʨ�U�덉�@��Pd̋>�p��d���5��Ӏ�t�ف~ehh7S '.���,�s�zQ�_[��*rG�D�z��A�[fRh��E�@ NF]
�K���ڵe15kI�J�*�e!$��k��*�,g�'�ˉX���Qm};�(���#FZ�6��
� 7���c&Ξ,���+̤�uo�R+�bN�I'���-�����g>����!Bu�d���LZH�_���ˌ���&8^z��8oCUtrr��O������y��玞<�r�����h����l�Sss��z�L�7oe��'�|���  }C=�dr�/~��Q��7�5���N}��	�0
$��,�##.FST��l8r�,���t,�1�O|�w߾54g�h,�=V��&�Kn	�A�n?6,|�������ҳ��,p��77�L��4�02���� �2��Z���[��*���Pa�
��Y����&0C��I��F�W��W�R���Z�`c���H���Z-��r�8~���3����N��4=^��B��?��_����m�nk�����T �M��" ]�����s�?���{�d��?��]�YZJ��gO��kX�a�/�Y�/Mė&G�n�~K(�������S��8�ꁶ��et�fĪ1�H+�^�X�3��}*�:�)�K8r������L�������A�N�E�"�/��X�"ʬT"�m��_C]F{b'� �$#.��n;jm�	�B���f'V�%��f��D��ϋ*U�eU��٩q�[[�U�ڜ��qh '$���W�\�:λd��x�.`)²�k�E��p��ߺ9�Ա�5���"�!�U�:a���믿2��y�����Z��8y�p�x�=_��WC!1��Ú�/��yt�8AX�r�	�ī &�pOmo�g�y��'>�޼y��w�㙧;���Ȩ��V*�}~��={w�3�>6V��o>��+�����aB��P��T׮�;���5f��2=<��bj�-�-��)5�����0�W��NO��*�L=�

DZ��&�JA��U�ㅕr��{��^;77�N� �R¥.dɘ25kQ���	���*�6��m~����,PsB��*؜�5�ܸJe/J \� ���J�^/m`k:W���0}���*�t�I����YT��lʻ�;�3�l}�C\"Ñ�/'�v��G��W�����p���b$���6B��%��~n2�]�GQ?B���`x�Zp9��o��>v�'��^�Ӂ{�,��!$ӻ��3Ο����~z���=T,�b=}����J� ��^*�Ӝp���h����ʤ�ȅ57��[l[yQ9P�B���2.��������)|u��-"�+�%�R�!9�Q$o3�����!4�� �@i�
��0-'�����g�
\����K4�e-כ=����@);�������
�3jb��m����Fϣe��p%��L��L�xz�"#�P�ܯ-�+úgP�fC1_ϥ���������;wt�KEn=<�0����v�*���RV�@U.�-w�e����&E�����O�p���P���{�èxVj	��ds,�m�>�����~��r5��?�%)�!|1v�ME�	�X�z�[��*��|U�i[���~2s��0&%��òF!���C�=��"<˺��'��eU��T���d�W=X��#�y1*��5-Z����3N/#h��K���"B~�l~E��������ZN�]��:�I���6�D;rhti�agU�* �ס:7�&k��:��w�_a;�FY�$��ܗ��y���r��hGp8���a��{���%�[�ٸAl�K�G�'䍬.��	����(KO� V�S��#���_}k�蠽�m�j�M͐��ҹs�WcV��������\W�@��.�"j�.�%�7
�[c)Yڦ��a\��j�A6HU�]e�u���9B��P���9Z6�}(t�ĎF��:�]�F���H����x�W���Hj{N�,��xE� � Q�Yw��Ɩ�[I����[��S��JQȲ�Ɇ$�nj���pm_p����1-�J\�a��xK�R[����+Պ��G���c)���Ȳ�i��t���sTBl�<jr�\����!��iʍ{S���v����������b��W��    IDAT��iT
�.W8�����P:=�ҳǏfЏ�DC�b���D�` ���u�a�f/�lE|��4���l�U����_��L�
�'� ӫi�dhh�r[. !�8nw� O�^�)���в�V}�
�rʰ9���Hԫd�u��ҕ-�o..���ꆑ�=*!'yH4y��^�Ҳ=|�2�*Z���hU>Mn�(i;
D?�U���8�1�X�6����3G���XΞ����L.���l[U��|���Ǖ���S8H�so!�+O���)�L�>3��~9�"��@���Ȏ�/�b%_�`Lb�]���R�Q�`7;�wdQs�$+�^N����d(<`�J����ُCw�P��!|7��N愈�����'�,��c�//D@�5d����Y����W���~J�;�>�a�7�s�	Y���
�T�
�r>ę����aQ'�����dB��c��H���k*C5�Is�f�E��ɷ�U�@ ��'<V��IS�Zt�ER o�j�-�l����g�h��@9�~>$¨'U��ʥ���I٤�'b����y���_��W��B�X\5c>ĵ����0:�4lC�_̂~���Y~�|o��j���߬���;U�U�ʷ�/VD����v_�8�
�P(:8�yvfa||*�F�=�*F#=7;��XŝF��?�b
P-�v����RۏQ=��W��
��c9V��PΡ��=.�s�5�E!$��2�iW',>v}�%��577�����E^X��ݠA##LƱ��lbryn�%�҄03�ht�v0�	a�.�1*ļ�Q���{�&R|4����m�hm97jJ8�P`������Cӣ��'48�
�l.��-��Ç; �v2��,1h��\0h,3QO���4�].`Lvy�01�U�#����t�T���'�֩mMТ\���43��#�G�uQw�H�Ű`�	�j_�� ��ϣ�S�9J�R|�֝���A*(^�G76����|�g�\qTjg�m�2h�ƅQ�,K'�
�겘��NL�S�5]���Ҍ��a�'
_���'}��E��y�!VشE7v���ǟ�������`O��G�-&���[)��r���y`����}��e4$��`���K�պ���*�S�<��L�F`���[��ɤ�K�Y�h	�^�0i�a����u�ёt2�:�.W�m�u��T0�:�͝�S�̐����M�{���W��>�&�C<j(jɎD��&5uw���_6@np��;�!��%��N?�+��q>ԇq8��0�ڹPF�H�xWAHJ�����2�k��������y�_�G�����#��(���i�?����)�������Z�A]Y{l�|_S�̈́�9�C��`L͋S�g<�2S�m��T�'���|��B{ʔ�`m*�U1��8>ZO�ti�����GB��c2���u��v��9�����"z��Q��pBޅ�0k�m���#x��J�;r��F҅�xO�j��%�F����.f�fgM\iF�W"�e��Q_��s��\��������&��G��$r� d3بK1� I�C����� [l��2��/����'#�n���v¥��U9�;e�n[��JD�p�E9��nL�0�F��ďl�Qb�++�
�<X�Ws%4w�B��ՋJi���ˆ�J�x��6)�6ĺ��A���7��Np�S/�<b���Ȏz8���p׃yC��!��uqq#=�Q��d��>7mڴ}$V����ry�{m� M�� $�=��b�Z�:1;3[#�	��%h�m97j���F����B.�0?�W^!�-��>"J�������>U���Wj�7��\��Eh�簉�}	�����s�dBI20IJ^XSbF��Ȏuwr#�%� ڏqx���Z�e�17��[[|�Բ�r6K�]�����E$d妒�T��Kel��?`��~�+���(�R�.Vf���DЧ�A
�K�m۶�}�6Ll��Lğ��᧜[�C<J�����w8Be�ٗ^����.��VJnUҍ��̀-�
u �|!�,��Hi� ��pb͙��ȁ1#���>���ȇX�1���B�]�2�*a2��.��z��j2����s ���2��R��g�,�n!�6]���>�I�!i|L��Xp,���R���6�����}i�֭C������O���ӯ��������H#1��눺��W=mO
�i~C�Ɗ�Kj�F�@5����溦e5�!ǀ����dce�!��U��MI]�p�۲�5���Q�P�\N9��7�!��6�3��<t +����
.�'p%�t)���	�sw9�Q��d�f�X��S�b{#��hQ~t糕T*��_�s�i4׋����Us��n�8�!?�5�`I����3Yu���z궞L6�g��\�ٷ'�Ͼg�Ρm;ި�Ϥӕ�a߻��+���'?}�W��x�d!�q���xi�9}�*v��"$( +�0W"��	�I���C�V��r���IU;Ա�6�u�Er���Z=���l.�r���H!��26�=\�ϵ,�e:^"T:o�&�l4h;�
%O0���Ԋ[��<r���4_O%�sڲ|�qh��
$Z��j^܁L!;�pg���
,Ƨ��ݿ7��ĻL�(/I.��!����9��%ө���0�&ʣ���q��8��)��ѥ�k�N�o��o��S�V����v�[�_dDV�\b��|�7��T�l��uo�-`���W���b.�wsC\��{L��i
H/�0ԣ��R�N%8�	;��W��]�.i�7��A�u\B�pqƃ�-97f�����/~�����?11U(��i�<��޽w|�w���?�����3cF��G��$����(ά���X�Q�:�j\���R�R���p�2pr�r��
��&� ���mY�D�t�`)�|r�+^�dU;p�Q��5?�nj�,���^�$h��zâ[���B��7�8�_�H*�۱s�Ћ
2+��FU6��`	Y >e�;�6��mVpM��5RV9��J��873�H��nX�tIߠ��G(g��O~P�ધ�}����|�g>s�×<}����$�����T.���O��3�{����ѯ��{�ӣ��0l��U�T���݌_-�`�s�:�B�����ĸ�?3�g��?�w�	,��yR���X7��
��� �-����³s��=�J*����8	�-�i�x���9�5�sizbf���㯅�	y~jK_\�j�� /�]��;�7833Cx# J`Fg��^���0X��j��zYQ��5�q��4IV"�^,�2����ɜ^�d�t�u�v]r�#�V�6���j�$��DX�Lm���ʗ�����������c�{���nݳe��׏�b|�I�>�v�}��_~���o�o�}y!	;���fd��=1\�� ��Μ{���*5{4ڇ�7�&���<�p-RnME�ۢ��d���SfR�fxvj8~�q��(N�=.)��� ���6�۱1�ۏ7p��SS��?b��\�E�IDP���g�
�[FF��R�(T?K�	]		c�S6��7KmMi
�r�F$_(q>��6j/�I����S��yt	R�l�C�(^sA�4;m��-���p�q襗'��n�z��{>5<�����K����cϏ���N�~����s�{�Xx�V� ������f�1G�z�/���2�N���5MV#�"_4��^cw�����څ�(�����T!3m�zLΒ�=����2�R�q%�
D���ܐO�ɶ��Y+�gf�\Db��(O��^q�^/�Ю�Tr\;É��bjdd�/�Xk��T��d��G際�5�%�%�j\�8p��Ni�1�⡧F?;ۑΣK4o���Pd�2-^���z��@�{�ܱ٩���=�}�'r@|�8���^��}������������gn.~��y�S�R(�u���.�I�k��A�=FN����Ġz7Z8���%4�r���*_j�#"�Ɓŉw�J�T�^2R�J���L���z���qd
0ٖ�$@��<�:b�man8���z�t�P.��N��w2�\��aU^'��z���, �<�aL�F��X��e��zE0VzH����@��!�����)�K�~���+m�J~���n�c�s��M��{���m9��"T�'�}����Ravf�,7_�z׶�O�?y2�I���`�5����˒h��zә4�n
Rh��W�TqlXB��7�O�p�1v��B�+��-Re�D �Lɺ��nO"<T����qJ�FEL�(�R��a��Ah��+�����#{�>$�P�,��g�+�9"/�tz8��Ė�c-�<G�c74��&���jŀWV-s��L]x�A�G�Z�r�6�:�.M��,Y�I:z<ξ�F$����j~��}���Ʉ�k�t._.���`t��so,�SK���֝��� B�\�w즧5U%-٘�n=y�̢��Q��Js����Ů:75(�����0._h�6W�0v\�A�.p2��Z "�ښ5ڲ�!1����>����/�S_f�L g��	Y8XUG{(��'�?�������v�	�d���@reGݪkz��mi�m��D1,m��^��PD�Yf�u���^?��5,<��z��S�=���
�p��üR,� �^�w�m,���?<$֬��r��6�9�!)��ٳ��_Y�`cg\��<�^9E��ʃ:�4��5�u���U���
;�����5J�^q����g9�S��j����cUa��O��+ԥ!b� 5��=�ؖ�A/�;$O�_*�7ۤR��`V��u[�o���M���GS	4�@%�]��Ź�r!�N`���W���Y@LԊ�JD��1��$�NL���ø��d2�]V#�2�㓦��~�S�g.��fJ���*��)4��r8�^/��No��s:r�U��١�ڪ�:��ѥU��\�c���ԗ{r`��s/'3C�#3���׽���{ �ߋn.E	���ȼ�e_���۶�R��t���P��>�	�慅m���Ǫa�J:2��J��Pac2/:\�y�5k�A�j�84�u/�7�E��+c�%3A���y�w�;�v)잂H�����܂��pm(�������86�E�
���<08��֌��]4�n�7t~F[�]�KF�Q���i�ސ����yt)g�*2�\���d����}�`>�¡�Wr��v:��d^;��ݛ�=�0�g	^ω�^n`0�30\��ffk��Q����4#O��04�dL$��M���Fy�a�6��\d�rǭ��j��t=�P47��7+�~T�S�(5+�}�f��c�T+�KF>WD*�p;�P'�@�S��h��y@f"0,���0��079�h,ɂ\�i��.eIv. �
��JT�e��U.�T1�. Y����2u8zaEu�`;�RdX��p��qL9�S+�⇎����_�9c�쿧\�>������g�#�R/e���jq��g��_}����H��'~}�g����j�P+g�iX�T�D9+��m2\�1V�V�8�Fp����>K���%S���~�"�%cԠ-�Dg��:"�>_0���3�i�Hd*���C�pwww�;����'��v�=�AWB`�"�7y�q^��k�Oo���B������f�4O&��/�m�Xt�����La�X����6#�ƺ�Zw������>s�/؍ڙQ+�-<
O��L6�/.����n��>���?z�7����`8�9Q��pQ�"��]1�:X)�ĕr̈L���N����S�a�S��-��ԅ��*�H�%Hql�`LR�mL��vy&����fWO��H���&�9�G��P��0(f�`��bܾXԂD<������s��>VKҤr����+0,�R>� �i�L�s�l� �i����/3{�ѥp+�nANנ$��b�-t��ķ�����ٵg����e������^�
���b>��?�F��3�艓��������36_�ZI�X�r��f����������n_�l6u1�<����
Ejn� 8~*t(�t��{�Y>_y�h���P�t�Ybo����b�놀�y<>�P`;��*0�E�_[
L0�	J�;q ��:��@�r�|\�`��ҩ�1s!��Q5�p�%��<��<z���j�V¯��1l�|���_|i�������ݣ�Xp4X^^J:���~����n���#�~������ሸ|�����xʴ��"�D� �*����&�[�,��݅�1�j

G�"){hSrs�"]�37����dKa'< 9C �]+���:��G�������d�r�JuS����F�8�sx�O&3�9�;q�e�+A���CԴ;X륪ڭ�Z�/��A�ǋ`]�̓x�!�D�A��u�N�2:�.����B�`p)!޴!a�X����ܾ07����?���>���|�;C8@�9
�>>���}���~��	�Jx��]�'0���.�j^Lv�`�K*�)�e��܀#׷")q�qWȬo�����ZjQ��R)H�J��`*�r��oؤX,	��{������,r��R��<�b�N�%Wb�"��������(�i��\�	Vx��^��D��)�u�]��f!�N�,�JP�|�A�Σ˒P�n,Vʜ^��&��^6\iq�lKD"����y��\/��|�����Q�ݷ4]�:�{��_�*�o2\uO@\n=�tʍ��G��.<��p8],x�á�=�c����O�H�\����S��ds3V�5=�)Rt���2[%��D�4}
@��h�(n����>�ЮE��I��D��q"��`"����V�&K����z{���z�[x�ꦲ��d�y�Q��8=F���[v�9�Ci��`��D�9�y�X��?͸���re"V�Z��u�,��z��U/��f0'���[���D/�T���ea;����G�8��&ytq(� u�HG�J[�C�G�����e.2k�m`OxA.W�f�~Ǉ��]/J(K<�~���H���Je�$�HU�i#�.V�bl���X������ g5�7���#������~����vl��YC���r��G/�m��:�t%�,�9�l7u�o�jwo�<���RW�lY�-/�n	uO9-���.����w��I��'c�\-�^����\t�ñX4�ŻW�a�-�S]斫��wcL�֋v!Ϫ�VT�U�K�77I��i+��`�v��w޹�R� ���Z�]rGK��|�v��_{�5�I��6rB�p�p�z[�jnL�W8q�۳��=\�tu��)���U�G�¦��#t��W��4��y��J{Yix����Ȉǋ���c,�]e|��I�B�� (:��$t��i��`]����
X��_g��j�����,ڣ�Z�0��W���������<J;	D2��\����N`��n'�w"�E���; J��S�]�����S�Y5�f]�*�,p}�����<�D!	��#k)^bT�g3�r%[(a?,�{¡�tV�>:q��t`A+�I�J)���&�r|h:O�#9�,���_ߘ���z�C��J@���]|�:�ۀ/���NWˈ�ATr���R��.3��Ꜿ�����D��z��]�/�.]��*e�:�.��_9��a���5.˘B�%�]nO ���Nɋ1<�s5e�m�9~��6�l��Tˡ�3��Vt�v�|�t��������iF�O���G�X�Ƭ׳m�fR���l^1��2�ڍ�� ����<07��qI�f������v��lt{6���ԪIhw;�.�"rF�'Hleg؁)A�d�^���If�g�܎\<��8xs����6�˹���a��)T�-��j|}u����	+0j7���ϛ�gկ7�n�߯Xvb(E�׈E��x���P0�+��
�R��0UsBl���%.���!-�R㦹���n5>���V�o%�F�g��o��k��6�;����Rɩ��Њ &x�V���-ಣC���\��ˉ��Y��p	��[�PΧ�V��ngo0R�f9���ᒝ+KpﵵE�=g7?�#�Q�~f�q��	�}�۶��#f�k�    IDAT��`��X(�s���E<gI~�Y���(���8�SR�����Y�U�Σ�

�F�a���� >@��R9[�1U�@�fu�]��y��d�*��j����[�J�\=�r�X)��._4>���T�i�B%��rNF ^v-�q��
m͏��F�����u�٢�v�[�Ӣ�K&u��J��U9L�F$����/���uNc�A���*��+�B��{���Z��~d��.�q%Bo01A���@l�]��^b�[槜K|ґ���ת�v�cU�U�U�V�0���e�P�L��[@��8�E�I� �C�4�Ѐ��[D�Նh��"���R-������3�]*�$�+�������s���|4�;pϞ/����^�������g��g^|erv�\��kw���C����{��N��xXt�f��r����0#N_�b؏�8�_���aoec�X��k�b>����` �#,|��7� պ�p'��������+��:{�yti��Z��˪�,ʹƨ"���=�\5�\0jK�G������}}��B�Zź���C�;#}�G9_(%���{��2ʎr���=K+p��]��s��Ϯ��6�#}1��-�3������β�:�/ݗS��<Y3��"�H!�d��6�������������o��cm�q`1&��#���GH3M�3=ӹ_�7���O��7==�D���~3�ﻡnթS�N����n�V�@�^�Q�zCb�!�[Zp�n��鞞����d2.��%�X}y��ق�����Ϲ�@.Q�xt�%(�C2"4�8 a;�#��T�>u�k?��7����#α]�?�/��׿��׿���n��>����NM�g�*���^��*�������ռ�,��y�?�~v�o��t�[��>�絊N!'G|��Soq�A\)����Y���K�߫�o6�8ۊ=�w	�G���:��\�_*����yh��\��T�Cϕ��U=A��D�VDk�'�C�4���^rKV7ͫ.[��Ʒ��F��H8[@Z���k���h޼��n��o����O|}��Q"�{�E��#��s�+�x~B�t�G<C��-v�,��� >l-Ur�n$b���$Őȕ�A=����� ��nu{3�?i��s�J!��1D��^�1��w�,������[��ɉ�w��_{2��KV��u�R�B����}뇱�C�\w�����
S�O���F�0��IN�j��_���Uq��/O+��Z^�uy���Tezܯk7\�����5�6ږD����B��zp���ұmL�R�$>�G�a'�I=PI�0���3�e�jImy����F.��gSG����'�Mq�6��iI��yQ@�$k-3o��ҍ7��"�?�����G�����ݖ��}��P��I���]_ٽ�t2�j���n���O<��a�Kd��i���d�
٥�K���Nť���|��vj�sn{ڭj�x�
���L��m�䒁�S�X�v�������ք��N�H�/
.G�Ü�>��@���K��*��v�罸\��T���=G~>�en�ɥr�ؖXn�0���U���u��xI"�;ڕ����[W�O�Vy5]����u��t���\8�Ɏ��/~񕣣��GN`�ac�4��9��f<w!О��N�-��R������G��]����x1���X8G?Q�t��e�"�uv�X\�s�C.	�v�����hY�I_ϟ\��6&0	$�Д�7��n��hW��.�Ѧ�9�߼rs�֌/^� g�����7��a�DD��	�0��G����e7������T��;߲edd����IV��@_�et� ��d���m;$�q:��}���^���¯N�թ���w��R��TO���/�@*"'l�)�8�:�!S���x�2�&�f�R��+t:�XK_(�u��1��]Z	��Ƽ�w�z��Z�R�����T'�o��M�����Ko �AhK�y�:#jZ�!Ǻ�D�d�-[m<\$G�*�rU)5�*L�c'���]d�J�#�%Zq�-����v��I���䋹Z�0�JD4��X�u�6�P#�f��x"u���'O !����j�i;s&/�E�F�[���E�p�_d�K2��	�Jx��ޣ�
����a�E�E�
q��� �s�4��;��.��=�{���SQ�����s���)�ӛ����|AoP�4_��d:���&G�@ȮT�\�����paR��R�#�?�X2�J�u���=�`e��#ӝ�"��Ȋ?k��I���\_��\xC�UDB}��]=]� �n�>�uC����¬^F�I�C,�#.=��0���f
1]ь��9���s�=�/,?��O�x@����Q��$�ʗK>=L8�r�(�k�p`�pS��>O0��3?z`|�x���P,���u��A�p2���������.�3��<]���[���!�#�"��#]|Io��Ze����')�-!��J�l�0Y?yj�c�$�%sEp�d�?�/(����ٺ��4p��%ČM�����[���4Q�ejO�=�+�C�65�+'O�Y�/Z���1?��Dl��wx�}�
+�w;5���p(�Lw�ٖS╲�g�6LO�`&A��="l��E�lq@�mD���B�z���"���mZ�a&��b��ǟ�(<[��%�x#xȥd�×L��a3}Z,� ���}����}�x��/����w�}x��>��������B��0=<=ur��?0�_~�}�����=��Ï�nX�h,�{Ä�Sn��n
p�۔ ��l���������Ƕ?��w��aN�^'�a��o�cbq	^��$��ް>>44�y�f�+o4؏��]�
��<C��yI��<���O.��F�j�J�/��J�6*M��X�|�����}�;o�zi���#{��ڵ�n�2Mħrc'������ǻ�����~졇�
T�Ռ��w�~T�)Y)��������Js�@8�����Oݥi�ac[��F�]A/��f
�@ 88pC$a?�"X7�o����]@i��.��ୟ��6wy~ߺ �R�\b�&)M0q�^��'&�P�L>���/}��ˮZsɶ��n���k_T�c�Ȏ���e��t��x<���9�o<�ȣGp�d���x%U��5�%B����^�
���52:ܕ��[3��|M�+��9d�csMl`�Ǖh%���}�%��"�E�Z�s�=�lK��s�\vjϒ:v���.�{��m:E>����f�4|�$�D���c����������?�t�[��U�����T(mt�ڤ9���;��|�ɽӭ`�����լ�	{�>�ɥ,��s�Pi��nk��~vW���,;�k�p�TO�z���ɂ�o?���s/�TH�E
'�	�Fnrr��˯��}`ͪd8�TJ�#���q�-@*jS:r�?���w�؁�&�G���\qknZ}M>׾���y�]�o�ɕż�3���v���s��^���N�]����0���t��3�9w�����
n�:}�
��\�w�z����Y՜�lëG�B��G�c"2HE"Mo�Z,~�?9=��7�qõW:�0�� �$�a�s���t���nYNW_�P�>YϞv�zH�����O��X��!@~f?�쇈.�2�N�^/T*V�~]�.�yh�I�����a`E�p�
��`զ�1�
��D�/��m��|B9��K\��*��\z��6�?���G��I��Du��t�5�U��#�݃����=v��"o��u���|�l<��?��R�����S�\������Z��Zn}+�*����}��p<F�Z)�!+��0���eA!�.gȥ.ir��!>��G쇸�����N�����r@���B(�3���n� �b3J$�˙% �R��؜��dz�������Z�ۅ�'�����.VJ�C�&*�X����Lg����c����ݵ�����mV��ʯ��lÆI�Q��Å��[��i*_������[��S�!]&Tn��g����Z.�b*��������O.�-e��W����O\$��u?g����z z`����{5��i��v��`(��v��1�ehk:9x5KB���?�����\�Z&�L�ݬ���QaYD����%ޑ1��r239�Z2/a-;���o�ʛK� �A�3�Rt��LǺ�䒷\j��хn,?�ʨ��E�Cg�V�h���W#�@��}�Q-���d ��EO(
���|jfK�t:D�H��a��Zs�p,�Ǖk�'�/�{���Zhl����D�	��r����93�zI�Q����O����"L8Mv��(r��%}z��e� #�F�b�{���8��r��ю7.�$�	�D3tZ	�y��WOZpjl'�P�It���e��������N�91�7�&|���L�L�)I�a��J��L�F"���B�@{��$�=�����&"�r=��&q�옣'�I��OW�%�\�rIa��I#WXI �W�<��e|��'e�5/����[~r�v��y@R7e�P8���g�T.�`4��y�eu��D��x*n��iJ�_/�����M����'g�2�Z0+W_����4��##�s9۱�Uß�n� �w���%I:�o2Q�+G�D��ǹ����[J�������sO�>|��E^9r鮷��]r]oz@2����n��u�����īn�L_��
y�����U=4�����Xlh��{Nwe���n�鵚!_,Xk�ysң׉�D��d�3)�|��P�	{'WNz�Ӭ6�\��w�]yμ�g�����N��t}9�(u0|V�I����wz�܏^螺_�c]�xש\�����d,I8�S�F0�h�sD��8�Ғ�4�7m8L�\�L[Kė$�����������<�Ю��n�ʹ :�+n���l˭p�����3��Y��gx�1�lT�cZA�9�Ǥ���R�]���IHTr	y)�8�UPlj`�dO`ۦ_V@���I�E��9w1�<rٹvYJ�br��؞�N�"bx��Qm�}r�fej�i-
��t�Gī�Z�Tӣ�t��e($�u8L�:BQ��_���<������}��C>9>~��A<(���Hyj��"���Y�X�+����)'H��������y��Ձ�'����Ԗܯ(�:@ݍj$�MZ��/����T)W�fXk���]M���F���H*�aS�CѠ�a��4�*�$�D |��N�r��r��S{:տ��;��l]oY>0@��f�$j�c����kբ���/��>����k02��>��\�A�r�%z�����g�O.E.A��t6�*�eL�ȏ��NhZe�7��J\�����N�Ip�S���9595��kɮt�k 7Z.�D�	��>[[����J�ez׮�|ѵ�^�V�����Z��:������@1%��]�X�9�$�x~�f��?�\��L�����H�OO8l���@�D��|۪��{w����������N5�ǫ���ß��W���R�j�Xҵ`���@�?�G+�W �t0��fź�u7��߳vm� 0�0�1-W�����!Gs��}h�-�ͯ}��Dv�z*�3P�e��tm]����� ����t�E��(�EC�	o�Z�6Mc�E�_׫�x�V�oD�N>|�a�x2�w�57�]�����'?���S$�>U��$y=�a"�_!�ˌAK�\wz��&,��jO��Lb|I���az+E��>]Az�6⥓��U����M"�e<N����r�`a<���RBk�V�Ɗ��)�c ��z�q�5�?��o���7j���{��7�>=r
YȻz��WW*W]w�{��&�Y_�����"A	I�hy}f��|���<��ܱ�6�=�->p�i�-���+�z��T��<���k�ך̦5�:��gGd�d���J�Ń����W�1��0-8����z�q�m������z�_z�b��r�D[�Uũ��Ç����6o��w������GF*塹~,4	G�+�緥z'rىk�����c�GG�̺y���Hh��cT�E1��&8��y͆�4��p�H�s����]�+�%�(��]�����'���ޕ@\B�F��;F�}s�n�'�E�T�6U���ʯ����V*G��'�ڹ�ʫ.���|$��h!۩L7����K_��[���������'�:tj�D8�751	�jԭ����q�qR9!��
Sa>�9�g..������ډ,�!9�*w�λ��?;���'���N�\�렄R ��
�X��:�ȋ7nZ=�i4r���\�I�����C��ވD�����㤠��٠���n����r�m���.��
w���#��3o��x�rjs�G��%�l��%�����'��:���K��:TC9�a��F�eU�\���6�]n�إ7/�vˍ���d���zoHcp����ի%˜�����/���>u�X0z ��o�|�}ҩ1+�a!�Γ��o�Y�n],���E���E�e�G�#���&����Ĺ�p�$�@7�����ݘ/T���xq�/Ыϵ��ƑAh��yP��'�XG"�Į��E�ĺ�%�Z��eە�ֆ[���DCk�/���t�����HK|��i�І�W�<uǙ>������Z}�e���;�0�Z�P�]��Y��"�sml�c
�����W~�^i#F���d�J#�әN��TF�Ѵ������ �(I�Z�1!b�nPL*Q
c5�`/���{�<��W�s�g��>k��XJ9C.ϣ%�\�+Go�]aBD��p�61����.<��N��ǹ˷��53�E*zT7�v�J8�'7]|����ٿ3_����%�@���FY���*$se�ss��ʅ���!���������ݛ	�(���K��b�L�)v�nH`��>o�s׮]0��T
�X�	^=P��䕺�m�R�Щ�M@���'�͙\zX����p�4�e������ݟ�4�Mͮ'� ��Ih��F���aMKy�ˀ�j�X*�#�H�Z�h����"w��1[yr1pi����'��|����=�_4�j�epϰz0^�Vjf �����x��nڴ	��fنß`t��s��e�a����󀀐��K�B�d�-?���mʖH<�5�|'8.B8��,���X��9r��Tn�	���خ[= kI/BhnZ��cF��F���t�'J`���8�,]v{�����>ǟ�N����\b�9%g����x�4	y�z����LCH%"u�����{uI)�����s�\.Z���]��#�H���̳�'���)�����$� ����S'n�拆��Z�<���\q��[��J���Lj��{�~��.�ҳz���|G�:rh����ɮ��4O)j9CYVHLG�X�1.�s/L��m���_v�K��-�$e�v�����B}-r�1\_��t	%t�LtA�"r��s��O;��ܶ��Z�?O<�����ҧB��mc�C`�$���}�SW%�u�>	��ğx��]O���[׬^W>�{�큤��K̃�u�2�b�G^rï^t��}{N?�����D���(�5���0�g�� ��?����y�A��f�v�՗�ƻ~uӦեB>���S�Ѝ�-S��C���}������!h(S�L|{Еc�93���6��{c^���}��|����gHlYg�Ȣ ���2nd����-���ŚA\�H�� 迓����vox���v�U�n�S����?�Iױ�P��Ԓ��~����4'����>6��ٰ�"��f5p�vã�:`kvM��tO�N�u|4$a��ob|*OG�1�̞�r𻎰*�a?T�WAV��>O+��*�E�;$�K�I�K�!vl�#�Gʕ��H�P/3u���G�@��T��Ȯ��4[�F��)�E�ڲE@�@W,��&G��IR���&�lym�Գ�BR$��S�ZIU���XN�����|��UΕ͌BbJ!m��>����6�������ʀLc����&�1��g��3����2�g��/�hUg~%ڙ$��\    IDAT�D���f����!=}�w�fNB����i��Z��K�]]��(c��ѺD�|Q���&�#�/0=ݳ{�n�.���W���V��S��sO�K)���t��w��͟ǳ����6�XlGf�� Uw�AN8�i 	H.Ȧ���?s�p�ȟ����׏����VS�1���ɇw!G���UN��f�m�INژz��n<�cS&�4��� ��ZXk����_���U��7�۲�ʧ�|4����>�_3�~�\�~h�ڍ��#��?|�ѝ�7D6�#ÇJu-��5p�>qш���x�
31��h76�^���`1�	6�S��q6R&���R)��Et�1�w8qi%�B�d�T
�6��!�7,O~z<F!�	)�H����ԍ�x.<���XnB�n���0�L��a�#�1�����	WrnU_ψ�GQ'��e��*E����4���C��d�R��a�sP���@;���$C��]�$l�O�F�\�s�)���A5�K� ���ru�E�Fs��ó5.�/�c8K�$���z1 5��B8�*�
.!l�C+�dQ�A1�PL��h{:��TH���<�S�U��~�xSp�w��1�0i�}�U�O��y\����S��q̦�	F������2su���]~r�Ry�!a*$T�b{�I͉����}�;���ӿ���t�����U��1����T�nٙ�՚�G?�����Ï��ĚH4j#���?C3�VC�&����� 9�cّP���¡@K뺿�j���	J�	��4
 �8qS3Q�S��LL����k)�iY5Ǩ��~�W�����Y!O��5Um�vr��K�5�Bs6�~���`d�d������,q͖Df܄"xL�P�0���R�Kǰ��B)Q7tL�D���z��S\&8L�)��}pN������\Rϋ����J*.@�&M��(��g_?���3�g���g*����=��EQ̹��������i��[�W}�F3$���xN�TQ�^���^�����/9<]�+��z>+.�&;7	�'�_�f����~p�}oz�ׁ�M��D%W(���Lq��"�-ԑÅ �2�1�TsPx�K/�G��hOW~�y�j�������F��s6� ���l��ݻ�S������]�_,������I&�-N4�!̊4�l`�h2��MO�RC�N������$��%��+�e��6���gpP6	r)VnK^il��!�^y��/������f�Vbo��B�>��"	�F�����W�4n~^�*$^�n�8$�ac�����Z�H� ���EFø�ȣ�,:��r<3����Z�B@>(,� �	gp��;�=B�f��m�g�_�{�����Y�O����I�y��?�
MN_G�l�������K��3��`��:�	�0�vK���`�ĥXA2�d-��VD�/a3�`���g�-}a>>g��A&�Y�������sa�ȥ�K��V<�*O�s����u�6�2ЖY'����q�1�^!�����'��FG�=�e75��Bj�i�j���5�n��b��ǳF�G�:�i�gئ]'�O'��;O��q,�(K�"V���r�e��}{�Ӱp.L$�Y�m�cj�p�;?q|_yz�H���!8�y�(dU�Pq��R�)�2�h�l����*sAB'>�R�Oӕ)�g����2��D��;���o�<`�:Y6�p���X~�:�Nh�l�\!GV7�F��,�#��#�Jb�f��E��V��N�(�"l�ee� ��_�!������\�ǹ���Lu�t�>��nsF��>������38k���L����L7fReyS4�}u1'�5%��.��3]H�<Ӿ�m#� wɱ�H�ۄx���d�v�.�z�t"�.����p\]�tz~�G!/�XAׅ��h,{0��c{R�����������/�$�O��^5t�\���ҽ�N��g�@.!a`3<��!*5��`a]��`WD��x �)d͇{������Nwf�Q�xٛ����z��Ѭ�Qo� ��������zi�����vgc%�u:�n9��`I	�y%T�M��xè�xV��\�נ�5��P������z��l}H�f�UM~/B�T4Y.(�V�T����O���U*n�b�D�4%9������<�a$m˄\Yf�)����i�>�y:o�W���#&�B���p�9԰Ħva֐.���_m�-�g�ia�h���k�HKڅ�R� �k�_ܱ�"ӛU]�Up�|Q�v�Q�����W��}�:S��T=SXK�@i������h����ݙ�^=�n�MVa�U-M��E���w��FX�c0���˕pD���O-u9Y�������<���M87ٲ��x=��c{���A�я��U��qgfZ>m��(+j��%{Ŵ*4�����64_�Lyu�a5jF˫��ޠmXZpM��	�<���h|^'���p�ܰ[�(<�d��0�.�?��;��b�N�g�K˶���-���5���>4��gh��~�F��� 5�$,��5Tu5�\B6��®X�0��r$'��ꮖ����Uñ\��>92��o|k���ɛQ��kB~����x���0��U���4e?�:��@��i����Ɋ۶���J!�sȥ�ԑ�Ș;�V �5���, �22�2'm����n�4^V6���Kq����B�f�n)rJ�B`�0Y�%��9�(���"@�����ԋ�%��!p�勏M�k&@�*k�Wg%a��fz0\�����8�Pb�8�ܓ%}w�a�Z���("���E+�{�K���0��f����L��C~_:��[�'�6p���K�i>��|�ӄ��mիf��L���)�I�1j'�=9:��^��R$"�E&&&׬_u���J-Ȧ�:�< 	'�$�
*����ȟ�c9���5j��}���V��h��9GT�_���ݝ�?�ѝ�j�J��s�e{;ͼT�G���dx��ã�]?�n��ձ_�%�:�d����:� ��l�i6l��h�[VQk�%"����U�K�O���y����ń�pn|�-4�e]�����߯��p"�PA�qV�G�wnE�h���%!ͼ'�J�΋<F^뜅�L���G%�*!�nj<[��~ȸ�V��X�_�'n��G'��G�N��켳�֍�POP�I����)t�Z�-��L�SgZ����<�s�@�Ŏ�e�y]�e|2��1֩�Љ��~���rٿ�������FP��ƫ�Q���M�*�����BG�fH��dO�E��r��G7�����t͙X�6��2�X2���-��5�Z<'�u���c3�'RCXEx�J쉐�'S��8��B���_��44b]W+ڣ��:q��7�G��P0f��c6��Hȴ�H$
��h��0j�O�鳻�ؘ��*W��)�n5C�HK�X�#y �/�����ҡ�/�5� S�Ee�f2�,�I5[\ٳ��U�b8��H�I�&2 K�fJ�D����e�u�Wa�\��Mض`�D9���>��R'H�7o5�;���:,�4^r�aw�%�t�cц����@&��ܱ<�-%����,L�0�}A�Rn��0�ش��d>.���۸-Vke��KQ�s9MNy�� �[�9%��J�h}��X�gE�V+F$��٦�����0á`"�������6���{zz�1!�Uc8 ��.��rճ�//��r���X�K��\�k����Qd��~Id�`D�X�G�ݡp`pp��O~�{��A�/��G�3�.F~�g�'��9s�|���[��q����):�I,�� A��݈�G��@+�!-���P��4*�aփA,K%��S�z�{�'�L��)��iCJ^�Uģ"��L�}F ��#����ͯ~�S���c�N�6�AY/�q&��k�F]�XĒ]$��l'��:��U�M0���()|�r���HB?��J9��L:������?F��T&9�����j�h�9P����%�7����Ǜ�&�ih��:����|��E��[BmU�bMW�?�O�fW2�u�6;<�he2"�Xؒ���i�lh� ��Ӵ�(JɮX8T��/�1����*b�͌����X?x)��峎3}\D�s��J�a�QE^�zh�Z��)��yYi�{�5�Ӷo�<1������3�󣉳�Z�4iW'�!#�h�xD���5��Py�A�ߌ��R	��zX����y��d�'_����������n��rl-+`���X8�?1Q��w�Fjz����e��I�q�H1�b��y�Kق�?QɈ/��p�+���X$ĳ�r@|#�FFp�)�D��%�5�^�d�kdT	��<�`�HeA�dNia�O#ȥx_0YdZ���f��
��9�i�Njd|��c0S�촰�ԦG�m��fA.vÈ���(��N>�hZ�iԽ]�h�ר�U��Qo(���0<��rR�9���	�Y�{�	dE&�P=w��d�H(5�MK�%7�z����֭�?��g?���;�@Foe�#��@ ��X�d����ғ3o�I
L�:u���[_}������K?����u�c�w���P�F��ض�:���$1B4���Jj9$
����e6y֨�3]i �T�����o�uC�l�E�3mq����K�����Q����~�TB�]M�����B����ƕ�5f�A��{�1;u<�^}���}m&�E�Q�x�x@�|
����j�������i�+�d@y^��u��,se	�-�Qef�E"FQ|f;�y4���aX����]w���cG>���#��o��o�*ޫ	G "�}f��[�h�/@v����S�	?ah�T�J����I`ò� N�d�
��d�0%e��}a�m4�)�ݴf4!�07��	��C��0.��5m �YF�c�d�f�"Bu��.T�Z��yQ#ȯ�F�\��Q�i5��6�@Y\ܼ-�,��T�@V�1⽳�4ؼWD� �X���C�RE���J�,�i3�E��G��kW�N�+[�2i���PܖK��Qb�~�/t�8o�]����m��~?{̭[�"^��^�N2Q �_C�\y�ຠ������z4��Za|Z�6�-0 ��<��A��H��S���ډ�X&L}i4�U�Rް�:k���9+_JB1�̍���~����Z�[��%�{��`�K��Dp!F�@�n����_��WO�8����u9�m�
ǹծ�/�ȥ;X���isg�����/�+J!{0I�Ǵ��PO�j��&����?O�G�a�"
0��G1��\�f�<v�]�8�	]N4;ұQ!�Z�|v�V��N�L&b�|������ޝY�j5�d8�=u&:��+>H��C�q@i,DS�ݘ)���4��}�2�>�#>?9�1���˿|ۦMCG���׾9=u�TW-ô���8��Y�H"����q��7�E��u���A�jE{{��izR�.�sq����Rf/�S$]N0*��
����AN�zr������^8�k��@/�FA�)�N�R��a>��"���"��X��=�5��߽�{��޴��P�;z��0�E�:A�b�,��5IWi:�C+g2��Ng'�����'�}�����%!i�"�޾rv�-;����#��4Bdނ���T_�j�D���W �.�Ӡ�
�y�D�c��a6/�\qzr*�?�Gq �D��U:�.O��bB�t��"�K�#2�Q��Уy�~a�\*9P�
 ܱ�A\�j�'�SL�I��*.��N�}�-�J��~��@����w�1���gZϙ��T���=�B��#����c�`@/�r�Ұ����(m7ݲq�@Z�d>�;|8}����G&��G-z}kz�Q���f�Qf�#c��~[U��,�j����V��aֈ���7����y�р�;et���|��n{��W�ڹ�~06zȴ ��6�24Sk�th��~�u/��_yW�d������&��0Z�J�1kߐ��Z��W5��'�K�ܫ�z�9��A��>�waNi��%�;&s�F]���25 �EE�P���ݪ0^4L��Ⴧ��$$�xQ���R��z3�>�Ah$_�^!��c�N�j�baz��/�N]o������@+&����Y3����$���Y���7��7<��Q/�{��eONg�KW�)p?[�*r[p��"����?j��~��h��f٥����m�m������*8M�O�m��!��{�,K%�K�H�h� G���dQ�z�P��F���׳! �͡���!���ȇ��(��P �<���\���6ۼZQ���Q���e+�k4j�@�%�����eh���K+A?�e\-2z`}.���O�஧�~�R��KYȜr�?d±�d�'��+��2%a	����37=0j�Rv@f�@,� 3G��N��9/�Z!���P/1�=&��|�vIN��;y��S;w��F$�$DH�P��?���f2={8]�W�lOWN�3����Ž�p��,��.ڬ`[��=����z���3�ϝ��8v��C\V������h$R�	���@V,��-[������ �s;�jI�M����׽��W^%�ѭsY]�r�
N-]�	�⿿0���>t3�|T�.&������G���Oe�2H�(w(������Ӿ8���Ŵ�7�Qſx�@X�|1KĽ��jy�;�0��S��`r���zs��R� p�W�ӂϜ�E�FO@�w`L�@lj�n.W+�H�)�J�*�N}��E���OX�Y�;�u'0__�ϷY�{���ǡ.��hw�갯q�F�/��;o�{~���ĩ�"2��&�<���.�r��W_3����H�\�kXY�M�ĊX�$J�V�]���P:4,�����E�YȖ���`8�m��V���b6;��>"TR�lT�".0�������CZJ�醊e�ؖ�@��a����t�|�q�{R�V("��R���+	��ӕr�n6�WB�b)����!.�T[	U�"h%��c낽=μ/��!J	��1���Z٣B߱��SH�mQL��G�"�r̗�T�����?�V��i�Ѩ�iY����wUsgZ�,X:p���ۇ��Gnx�U������?�����7R�M@1�+?��;�#��5�d*�~4��Ll50��݆D����@�Ny)� ����_Izq.��������ʯ�����iF�
��G�L,Ax,+e#��h�H406q�c�+ì��?�y�E2�b�. �����ډ�v h�t��ۗmؓZ(��7oN�}/��w]jd�rx����Uo+Ҳ��}O~�꫟غm��n���?|�����>6��g�ʕ\�q�f�b��8��@oP�i6�1=j���f�A��`׬�-��"�F=���i����sYC��1L+�>��h{��k3�� F���s�֭"L֬� O$�OOjv=�N��j�K����14$���,�~B1�W�ad�$�Z6U�,V�Wl}����Q�Y+�{�1]�t�A�NE��>Z��\�##��"Ԗ���F�V0	�6��������w��}�O�~rס���F�G�a(� �(�D�}�F�l�\��5^OupU�m�I��6�ߖ�/kj�	� ���F�8
��X�q��%�s�Ԩ���b��d��=22Ft�d<����`]mv��u�%��K_|����N�)L�B�x8`}l5ekp�b����+TD�{����8$��믻4�d*o���ދ&��`��6C�
�%�7z�X
)��(���"�B�ث���%���Ɲ�󚱼?I�� ���W:}E�,�t��A�s����k�B����CȮ��DUz�Sj��[A�?�����a�]��/��@��3����j#Na�Q��"�6��ц��J��aL�#��j�Z�ɏ������E�N2��t|�Y~�R,{�)"e/��0��Y�X�Q����W��57b���#����ɉ��/[�j�Ԏ��=26>��^v�moy�ٲ����)�2��a�D��-�(���h�JɎ�@e�$���    IDAT���R(�	�b0J�`�;�bH�2�~T0�*��5F
oJL}�!�`�LD����I�	۪�����
&�Z�D���R�^��}i͓�q�2�@� 2@Ϳ�ܶ���}qOF;}r�;��棞G�+�>�<�T�WS��0#e�����M7��;��"�>�����Ŗs��ɮ�قO��B������^"�uwezz��a�Ph�ͧ>���~Of^q��S�cGG>�+� �[�v���6o�R-���݋Ƌ�6��<��{����v��k�nݺ5ED�B�Z�"���C�yϯ]y�EA�+m���N&�%��Ii�:&���T0��E��C��bf��!:��!�NN���-!;9�6�
:@\"��E
J���j.-�?W.��md�)1+s)\?�z>��m�'ؑ,�(���"���%�r饴M�4�� d�9c �z���011�f��&��2q!���x�<Y�U���4��^�v]��D�ǶF�Y3�=��CO�ꎫ��� �J���O��"�n�	����[���M��v����=�ǧ�[.��տ������HR�������(��x�p�e���#?|
�A�Z3i��
-f��b+�D�P�T"�J]FwwW�@W�X��p���+�oW�M��U�&d6�H�z4��Їm�9���+JJs�Y��!�L�Y��z}:!1X"al�q�a�1�Y�0!�j:)������Fwwxj�8�8"��ނ��S��{�n�>/Wa����q�#G������v���ӓ5�
�����/U��)]��8�%�A4м�X"���S��wϞ}{c��σkN\b��.����O���	H0d�]�]V��L��-�0j�(G�J$�r��t��cG�_��[_t�E��l��b9<[4
J���k���Hd�ݳ�ȟ��_��&�A|�0#�3��>D-���_���Q���aY�Z�7���;�J^�q��ڂ.�5K����\��� ���
��D��YG%��3Bu$ȡ"��<1u�X�2/��>��N�Y%�QW8Q�#���&O�4f�<���!�t'	����x��X,V�9�jcllƚ^bs������"�H�+$Y�we~Zt.�yi����3���X�[׭���]����c�=}�n}��Z�m�Y��**�������=�=�ӧ��p"���UG�f�>~�zо���H9BGܣpV�h6cAb�[Z�Z���`�Z���j�V9�bq}� �=$���{���A/��	��b��r�X5�(��x��l�+Ӿ���3~٣5���gS9+�] l�i&�]���]��#����u�E�6]���c2J*u�z �r!pi���X4Ƅ�>�f�V�����0M�͞X<MĦ�vKpU�_�+�u�d9�&1��	X��ʁ�G	�D����Ox<���$�5b�������_��!��ɮ�6[v����,6
��E�鑑S#�:VO��3#�)�UfT}g][�o*�59y�K_��c��)�O�|s]f-S�SCo�W�X�n޺D\����/R�Z�=@�O$�b�,*"��\�#�gh!3:|��4 RWsY�HQ�٣��,�(��]�Q�����f��&��c&H)���k�?�D�Ha�!?���+����U!5�Ù������(�%�c�~�jժ��~�T�j���rȥ�}�1v��Ź�;C�K/�0�O��GJ���ZkS���G��2�v0F���o��F�G��t���p�֓ǳ��NL��H�^�I�R�٣�)�;-ķ���ܹ�������{�P��>u�@���4��o~�F��b����ۇ�h��qB�Oe�z����?����|T4i�d�|�1�@�w_/M������M�s&R��,`e}c�	s���|��]+����5=�f�qQ&���:SA�lYN،�3�lA$�G���( �*�h,O��E�Q�\NJ����5�e9���M� ���#��C܉)�Y�{#�f�gr�%W^z�@�<��496�y\�u��`��z8�җl��%/é��wl������ @��!1v�h�<�)��h8b"�9�ۏ-|"a�P4�ۻ���{3Z��</<��u�K����>$����%B�z��E�#|�j��s6]e�^X���UV<�>�xő��X��\��;�y֍9p>�z�˳�w��x���Ay��D�}����,�I��8����@��	M�Q��o��>6|��Cf3��?��K�>�=��a��d�H����F} �tl|��gw�B�]�"<3:5w��=��&Ih�=FI�+F��47�\���T=Ѵ�[�n�.�x��!��@��z�?M�m
G���,��]=@\O��%�93{�B2��L��m7�@��s�r����V@J2�jF��Z���:����X�]�~l�L1{�h9/!�Y�FǊNs����4I�c���uG�P%��R���|w)�;�x�p$�\0�5�-�a���8�̲��>��ˌ�� ��F!W���ǲՏ��H�@1B�tTDqI�\5}�u�u��N�2=���ِ��+�����w�s���r�_����4[�*�c��چ@�#�k�����}
�/~yM._{����i�t"�WW��;0�{���Cв%�:�h*VPp	ì�OLm۶���� d,(�K�H<_ �7�7rn\0�2E[{��)���$I����=8$�d@"	Û,"�b��O�psq�Bݝ���_�T=m��s`Ac�R��Ž%��_Q~���"���PK�(K]���?�֧aa؀�Y}�Z1��ky�L>of������S�L�x2� �MT 6���طP��Ꮠ���C�x�e��Dxp�&�)��~�i��r65cl�8U-��D�%��V�����-�|Q-��	Pa�`�^a�A��0�≨bĨ{���*�.:N�N�_��n�nt�7�V�:~rdm��LW
�x,42|
� �-B]��8m`6�2�DP����{�V/gs���;S���f�8	o����֟�gǖ���ΚmN���&U�E�:Ar-N.�t����q�����Ya�E&�I��}Iͷ�_��7�D&#���a�믻���"�ǋS�B!k�ƄM,���H*��'��l�u�Ҫ�o��J�Ox��A�����R6�/J���F�(�xg	����r��i�zDXI��&٩�c��ކ���^��h�=H3E}z
3�p!���R�m֌r>۲m�Ƶ�z��"j,���
-��	w�U3v"-g���݋�8/�3h��(�}�߄\r;����jV�<0����-�KA0��*�p�522�0:i�~�M:ݞCguI��,�.�9��BC�!�|E,c���Ik�)���
���hBi�K���,�N�pp��7���#��o��o`���I|0�����l�RG<,��|�⢽���bً*�ٵ��a19#ͭ(ʽ9\�+�q!@�|>�=�?t�'��a+�ޛ޷�\+OL���}R�>�3���b�����6%��^4�'O���ޖ�����׿��
�*6e*�NJ��! �M �����}0����+_��`�y���Hֱ)�Ɉ�P�8��ܪ���e��5$��O���߱zuω#��N���c4>�Dg��A�-`ǜ_�W��/
4y��	�No�������&�ڽ���������W���Bxmȷ;�]:.|+[�f*��D�L&EY��I��r�Q+�}cc�w=�o��c���+b���T��Ԗ�K8�NOO�������
<emO�P�%D�kE�{jf�׌%���C���`,f�>�555������Ɩ�dEu��cP�8�Q�Y�>*�q_�,�-�Ǆ�80�ت��J���s`�-.�<{.�@r!� 7���:]����"Dv[v���K�
����lde�ㄍlUlW���LM�d��|��~���۞�y�/?��/}�;djX�f3��1waN��T^>�h����ƂPZ~r��B	�ǆ�^��d&�h�G�?�淾e��˵	�Z-=��+�]3��W"xe�J0�ٷ����^|��Ȍ�nY�c����@��ff�Ee���C�XZ�C"����e�����`��CaƤǀk�=��Go�h���"1�L4j��\����!#����CA�	�I6�d��V�i�v�䓀|�A�(��?'��Z ���Sh*FQ�W������ņ��&����G�DR;�R1��c����C{SD#1�Y�� ��A����b�F�	S
V����7�
�l�R,��)� ����oT(f�,@Lz�6���c`h��ќ�{$N��eW{z��Z�#C�5	�1�*�� &����X�x��
'P�x�R]_vz�7��Q���"H�*�Q�>ڽ����
���W2!���a��G�H�Z<��'O�<B��\����#�vޕs��{E�zv�]1�P�)���DK	�{�΂��-��Bh,t��K����]�^�f˅,���׆I�X$�<���#p o��$2�Dy�:�m�����*y7>��o|ë���֮z��-[/��1w.��b��>|̯��Q��NWw�^�v�V�3���;��"(���.�U�D'����/�W����ʞ���]q�k��l߳����G7]u�t�t��;cçw#-���^6~�t�������0՝��J£2rh���ꆻ�j-K\�0z�$���o��m_5�Z�v-kC�`<��V�J[wL/{����l���R��Ӛ���Ţ��z�DN��H'�xdx�X�8uц�Wl����Pg�P�S�̣ pZ~���_���Px�8���+�/�]���YEf���<�DčS�����u�]'O�"]�$rd��q	a�ĩ6M�1-�i��HQGw��-����*q���;�;�Xd�V��R{�<�O�lUz;� �m��f�2}��7�gU	��Qj�!��g�V���� �%!�0Ք��ݎ�&��\0���fC�@	�:-�rӠ��q��	���zM"�ƀl�Bcܟ�c���:���$�w�M��m�ʗRܥt�7�rA¸E�\[���ޛo�� U�Q٩��S.�U2w�v�}!�̽ڦ�s/Μ��`�'�Fd��sh�0�t��1�� # ��c8`k�s�Poϱ�H�5}��7���?��+��\(���f�N����$�Eg�������M�^+���>ł,��E�,�Ǐ���:璭laQ��$dw�� R��c���_�ˬ��W��_ݿ�������O��}\w�@ �jX�`���\~勴V��;�?��#����1b7FS-{�'R`(cO��Dԗ�db1���ݻ�_��O7ӵa�L�V���+���O9||݆ͫW���F�jͬ��D
�*��f}|���&�GB���u3}��pp��'��n��zׯ�����l�;EY����rM�7#}�d����J������h�ڣ��J\��P��\�VB1��)�{<h0�O�iMĎ=�0��h"r��Wſ�g��	eFK����5=OEM	</!뫄��iN�C������[�nM�R�g{�r�b!s�q7'Υ�}Y�#'��by�iT���j�J~���)�	�|Z�D�5[�)�qk	��g�E��h��;��S�GV�a���|H���5�bd�>5��]�ʳ^H's�\2zz�j��S�\�%񌡉"Ǹ���nU@;9/&�]�nF�[BL	���r
�PQ����*��1�IDxZ����\�#��D�E{̷�F�w�cD�F���4�pc8���X�8]/�e|[����_����kI,�!�����~�����&�z��S'��s��@3�B�H�
�H����̰��h1�������Հ������${.aU|�=��}�{����m�p�U��cwﻛ���$T����/��'��Ԓ��`�?}��>�x�l�kI��C_�읙?j8��'&��`
�92��/|��_�:���t��'���A�����_e���x|{8��$
Ŋl��\kA&ȯ��af�U���w����Q����c�X׭�܀!�H.�7��B,�b*�#�	�uLX�-�b`�]�vj~�5M�����q2f�3U1��X�5�����_LV�j���6	��%���kOtI榖�N�|x������j�����,�x��1�ҳ1��$۲h@*�s����;j��`gy�z�~[V���F����%����#�@��#��)ʉ�p	E��f,��'���@�t�aC��f�E��D�Gf�q��h�	��%��X�QN����?q�2��.�m���{���j�[d@qU�ɀ�-�D`ѳdq�s�J\�U-LD�L'� ���C�<N:qV�t�!pb�����i�
�a�t�X����a���0M���<A2D�oz���/ }G����}�ӟ��SO�fFc�z���C�lif�n
f��Q]a���P�����s��H�ǌ%�$긬�MO�g�4Vٽ��w����zѶ�[�����!��^o��]��k��J}�OG����{��x4\������<;3u��3��4�E+Uю50Ud��g�����tuخZ�ư�h�ر�^��W��8�J�S�v�������#�Ø5}D�I�
������g)* ����_��0!�`�X"�A6փ[��c�5��� (���(m$WȒHZ��˨�9�ۈ	�S����+!2Ws����:��[��!�@E��ʎ�%)&��H]��5�{��+�Y��"��9�삲�il��{����=v���ٯW*$��s�x�}�ĉ���;�9&u d&34SY�	p�T�~�Nl��a9�@�Y�1��m�Dn���S	��r�Uq#��˕b��J^��zOO;�������*�|�R��Bl�&DP�%5�V�����@��D��VD��W�I�A�?�<'\e+�ٙ(�gU~���̏{{�gX�(Pd�sg��=�*�a�*t�:����
r���eM|�,��p��ԫ�R˲Q�	�=M��%6�ƭ����7�]�E3a�<���'��&b�$S`%	B��QDeg@`�z���6j���J�^~r�d�M�,��[R���[��%F�A��FG���̷~��;�|ͫ^��UW ?��1/�J�Ç�>x�=�~��5#���*T��r	d�b�2�n��G7T��(�V�0����M/~�c��OL�����u�jsj|���_��?��W���{���_�����;L�b=#��yJdi�\�y�����W��bѹ���ן?5��'Rz�S���l����5~���Q����!��N�ض�%�ܘN��q�=�ٿ
�~�ݧ�3t�B��E\���"�q��x.��7��W���ѱ��w�=td�v@x���V��܅��5Qt8��2�,1�tؘ���}���ɓ�T(O�^��(@�+�?��4rN[�D�j��e覛�O3x��(o�qP�u�V)�tu�����y�������h�^/9>r�C�/ٲ�dz���NH��5�d&��b(&��j�0a\8g��H�'�i��O:|H»�0��Ĵ`4�VF��"�9��h���>�^�=G�D@�Ȏ�E��H�غ�iJ�EH3����Q��G$@�wt�����$D���S�^�% �!V,%�>�B���kv!���K�A6a|B��t�$�썠1�j���!sL�1K��=��?����&'��z�&���[^2�f�Q7�E\c�Pʨ�Zd[<���@iy����ٳ�GQ,�E�K8A_���O.���P"K$�Y��Z�MM�=���C=W�`b����O=����^��/[M;0�dR�>5��΃O>yrl��R�{ggWU&���k�ړTv		;T@�{Z\P�]��U��E�ݵ�G��N�8��3JϨ0�OE!�K��=�Jj_޾�o��9�U�����&�6]'�����s���9�����u�0�#�K�#��� M.�b6`bj�;p���`������    IDAT�BP��l9j�����e67�C�>���ݒ�GҐy����� �j!@WDK��TADlM'r���d3$�1�͉�oQ���"���
��[��� t���_��ug��������޷O�.�[e���&��XHۄBX�� ��_����n",�c�o;4H����]V'�
��0�5���q(9D2����x,G����dRط��X͘�|���\���Ղ"5W�΅KīA�$��t�uX&�U�Yb��7m� ?Ab%���">�QBD�ҕ��	�K�'���|��?�y0G'pr,�v�ݼ�F
�5�����cӦ�3����$v,1B���<tdׁC;���� �9�YD�)я�qT��h��Zl���C�����5�#� 1i� ��P$�P ��SẠ�1$5$*ƲN��q��sEߣ�AAK�]c��N8<,K��6 ?�
�.��ZP��N�m�A]�ʎ�.�����R��t�`��������vݵ�6*�!�*Ş��|xK_�R�0�=���X��+;��@A^2l��-p�C��GF{z;A��D�9�38��R�d%�H�TI%� ��+��+���
���25Ac]m�p���=��_�Nf(B\�k>$�ڌ��D㩸$.4T�89�;ԯ^�d,��*,A������v�c ����6]����X��!I��x���[�Z�ȋ0�56��64��H����8[��i�$S1($�E ��)��e�FR{��'E�s|r��=6{�dJ�X�T�ڽ�#�^9��"z`K���$_�ȁ��FF��񬷔��Æ�|Nҟեô]=±:9:e2g�D�I�q|��'�6�@�9��cՊشʰ1�T��󺖙^A�KQ�i�Q��qƷK 8��8hxh4�E�yY������+5SgגTj����O�8�,�R�Na��� h^���0�M��KN?�LP'�	�+쥔 ��DMd'7��XVN��!�B��=f�QL���V/�H�[�#���¶�"P��o!}$��{XD�$�;kަ%h�Z^������+��=P�����[^?Y�3C$P��Kf/i�dQ��>_��ܵ{2�#^-��Zyۧn}����8 >�h���w�z�Z��X�-��-q�ax�b�p�e/�t�����ݻ�B�B�c�!�D�5�Y���z�s�Ĺb�9E%56�GF
�A�Tt�~xG�j�g�RK.�)�7.�eռ�����C�R�K�I��g%o����P\a�1����d�8�V�d���7�X)+cn�f��nbn�c�`��kN��@:H���#3�Nl\�/!�"�'��6�*a�hvKH�̙��X���f�u�D��ʆ>��~�+>�dDC���)2��ي/qQ,�JP��b&�e��8��o.8k�[6<�hlh�H�¸9���X����Ӷs|���H�f��+�c	�"����z���N� #��i=�v��@U��~���&W(%��ye��)pf�$Ǚ���L3�b�h��\N��=.����S��_p1K�m#�̌�`"�
�'V:�\�|%�$��qf;�qLv�f,*�� p�E�I�'@���2ۖ������S�L*p������*UB��J�X���j�=����^p��
�����IZ�x��V�)��Y��\a��ႏ`�XD�\ SHdx{�`=2:59�=�4^p��9{"d�L��m�Tk�W��B�C�9� �_��&b��*�]�.��Ӕ��K�g�����Y���Ofk�tm���+�8��>زTAr�d$�7�@Х9����Q'|��"a�D_'�
�C�I�r
�nN�:���h�fV9���SK�Y���c����DBr�r�E��KL��L�d �J�!�I�� R%(%�ꀏt�	�ݣ��J�(�uv���E�!���dpAd�\0��*���1�3�h,�a����7pl'F��ߔ0�`nUk9�H�j�p�T�~�r6��NM��G���._�K��.w<I@ "2 �Ӹ���ь�5�N��D,�t$b ��E����	L����p"��D�YM�՞K��N��A��B.���	���]ٜ5Ԟƨ���a��4�=PPCĎE�^'e�^[C��!��?���+������A��ae�㋙a�� �"�?�Q8�'h9�#�MI�
�l���C��V[�c�f'�l�3�^�RQ�H��E��j���Nn}��w�h�I�p�ut|��r�b;m��R��2P�evK�J�
Ҽ� �Q�����^�*@�eu�E��+�j�P�#/����ʖ���˖-�&��Z�\��ػ��u�N �G��+-�+�T�L��q�;w��gdxlH�O%f����Rrc�N7�-MV�� WU�E�7�(��uY>��^Q��[C���$<��+{��CԪ�6$&�x�C���W�z��:�<2�XҸ\�ǎ�����IQ�3�Ej,xS���q"B�=��Y6�X���j9�W㉂��T�"��;���������M>�������|=˒#޼z͚����bmq{����+V,��:v�O�9t`/���곷�4
�4�5A��>^4 �O_RS��pY��i,=!V�� ����c�)�=��;n��T&��oUw�l�*�&!0 �(l1ڐeV�){'����F�d#ڵ��ѱ�뮻�#OED��wg2Q���|�T*ςI��aX�ׇ�A�/�M���xl"z*.�S�8i��31�L
	�#N��K��ډ��bX�K�bn_O[��U��a�e��0��C���r,C�zQ��z���ԩѥ�"�Υ���X�hl�1�/V�Yh�^L�!E18�]M_�C�u'H�H ���7W*�Z��r��-���������BVf�&�q����p��Y�NFF`(���~��M�uLND��1�&F�k�P.�Bs��梖���]� T�Jo� H��h�l.~[�<G��h��w;ۣc*c���T#XZJ�Q�	�F�B�
n��q"'���*�N��r��ys��X�q"�,_��-�݀!���D���N ǵ,/�T4�Ȗ9�J��y��|��^N�$�J���숈��F[sӜ4�eUt��uxyN���/��?�k��x,��{��u
 G)���A��E��"���Ʌ�"Q��v��� ;���'zh���ç��T����%�K~��TkΑ����뢱DAb	��+Mt'����]���R.����N;�P�v���[�{����.������Ԕ4��eqxZ�/������[^��O΃�=sӺ�����8b�"� _0r
]�� t�rt��ꗾ��1I	����l ,,ٽk�L(��a�c�� ~g�.}>��%]GF�n&����	_��7�Ld���֬>���Xv�l���N�����k�[��4��1009&ǧ\��h"���0xs�*T�4�G�b�ԪQ�����P�-����eua�$�k3�1K�C�L��P��0:�g�R���!�2�10�7Z�I��k2��ߗ^�i���P~; �C;������/���s��
�� �hX>x&� ���v�F,S���� s�ZE�"G�d�=�/N�!��>1�<t`����}��W%��X�pH6q��ܺ�"�j�EFKٝN�8 SnA	E(�D(��T��O�]K��=+��s��a�&����G�$bj��ٟL��EzӪ4�����|Z=�r���	Ѣ.��缑?sn-ti�~T�s�`PF󞟾�oOb����X$s��u�1N
�kR=?5GC ��y�:��"�`��;t%C����4������۾���]����p�wI�[w|y���z���|��=)B��ln�����M���d	fsP����]�(�����X��.u!:|���2C�6'2`R� �> ��u��A?�r�R��V0��(d4�������ΐ*�[�	���%������ ���9� S��z��r����<Jf}��t-��	�-=4�y䡇��W�fr-FJ�I�|{�ȓOnɦ'^޳c��H^��#���J-�F�j���M�����:C(L_|q:;a�b�w��ɩ����5��p�On} �k�j�R�LC��� �Q!����|����/��P�1xt���z���OQ��XN����W�hQ�]�d�י矉!iևG'�>���C�v+�1�*hZ����`�����"g�K��N+�c�H,o��iko#�>>CC�x�AM29�P_ȇ�f=��b�X�1у�6i�IN!�ۅ�\�����W*�=�If<A�D �=T%j��O�0���.�����N�Q_��$���7�%mw�9I>��>�q�!�&15!�A]f��~���5�>�]���i�~e��;Mc򕂓H�����J&���޽��d��zĚٻ��B�S��rVa�Oɑ�m(5y54%ݔ��T�d!^�_�A)�G�=���;���>?�*������#�/��'���V�_mV1� S,T��-�ZVE�O #'RGa_]��
�"�B!�@�]�LX�V��3��������m��N΂�h$�M�MƞkL4
�N�O���
*������jF���"�A�KA��2�-t.~B��e�E��yqY�T��Y��������hx��l$:�I���S�O~��w�E��b^e�h���,��HA�#C��o�L��2��L��KG�^.���"�,���~���SM9 A	�mH2���/E�1w9�|��~���C�Tܿ�E~�(�,��9���s��Q��B+i���s·>�w���S���&w�܇�X��pD� j��D��f�/P:q9a����-1�?r8��O}b�s[-6�5��C=#�#��%���Y���B�VD]blL9p@1�LM�"@��j�YJ�^@T&�iZ�'>q��>�~d�8��l������D�� N���F���O�J8�q�"#�b5j{��6OɋU~n���7���!>抳<sHU�D��s����	Dg��CN��\�cT��IYy�ʏF�M(N�&��V.f�-�+����J-cs�t�!Z�*�+������X���F�6a�(��hם�[S������U��ί\yv��kS�{}��u�W�1��X����P�;ӝw|�ɧ��r�=��p�''���i�1�=���&Y~����t�Bl�E�O� ���n&���x�(!�8��ʡ�T�v7b�\)�N�=���\�W򧄜½��ѳI�U�!�8�L�vCњq2�!g���V!ad"��x��X)�v	�.�GPd���m0���37�q�Ȁ����V���0KZ�4�8KT^�X�rPI����`]:��zȎT`z�fAĆt�Z3�q��P��l�o�Z�l�ˍ���G��T��*AY�E(oa�*4J�T���y�wO��;S���Z/���r�:��o���F�'�(pÊ�ᇟ0ۺ �6��1Ю1{��O�ջ騲F]2.Y��WI	�n,�x��� �zp�΃��sƜM4�><L�������tP&M)9�s8��]mł1/�����5�6�-@��� ���
��g�	E�S�D�"��6	�@W��H��d�!q+Ȱ���^�1L$#�|�D�N�ԛH�N��ޯ��?sT�^�rӬ��2Gxd6�P���\�W�šf8ӏ�:��W?}�s��4��x�}�v��(
�Y�W�6)=��r�2Z_<E�Y���ա^�l`�17�&ANV	O9�E_gGw"��7�jv����ů��.�=��1�Ϳr���ۈ�O(���%4	qo�ZBXW�����([��[jX�l�h]�E�Q8Q�Z.�&r���8|���`��Sig��/i)s�Jz]8�r!��N�Q��H"�}|���%6Ie!iq*cj�~?*P�U1��VȖi���(�D�}���-�Ã۶m߼�ʏ|�^��1�xe�02�B(ԅ��e	���'�'N»+��l�c���2h�tW�;��c�?{� ��G���Ϯ}�-�ъ I
@н� ��:�*nw�141:`�@�4�09{�n��z�5��}���p�2�����-����'�m��<�Q�Jh�5��e�5��)�RIb��"�x$j��A@�%���޶�)���L%�^p�������w��<��-��탉�D)������p�>���7���5�ox���868�fW�$����K�,G��d�>��]J=iE��b�"E'P�IU�;��*\=L�	���y`�Kze�"���f�����b/�����0Y�q]�����\��[�j���U����
ĈL6�����Q�{h-J\O�9GP˜+������ d5)����������b8�ᛙ#�]�g��:�Tc�W��	�R�o�#t C�%_͌��\�����ޱv�W�q3p �U8�&'����5�Z�3ڜAa�s, E�/��K0�^�
*��*����HS/��S%%os�ӹ,�Vu5S�͕$�- �=��^E~�����۪���N�cW�G��㓤(`��3�,�h��y�uA�����d��ٴ*O2̙L9��g�L��e�լ�)
t�)�R���fh6�ĺC#g��K����p�w���֭[W�}�e��r8�k��qǮ�-���BU�XS�����%���a�0�($n���W}^��#bժ���\����;x�ޗ�>���ή�k�$xE��,���R`�v������Q�t��k����Lg��U��&�Rd�볓xd&���2��"Rt���r�M8���合W�F�q"ܬ�-
*���0�GG�o� �%ӡ$bp6C�=P�J��3{S�qї��]q�E��ٻw���x6o�a�a	�Ld�\za���������)��4��c	IZ5E�X ���	��G�xbV"�b�[Ȗ?H��ő�\���@��i���@� xfGf ���d�w���P�i0�u��x&�Z�T��3��iac��y�*G�Ð���}D�6犾�����e�64l��R
X���v����HZ�ґ�SW�]� RS�/ŐIT=F����]��H�����j�E�c�=K���w��tZ޷z��C۷�E@��s��$[r*�T���)�+ tb���݁i�6hZ }��SM��򜖁��ˇ�f�6Kt F�˝�d>��e�A�c��d4
A�����ċlD�EY���͛�Y:�@���W/z��]��xBd6���~�g�={S�����_|�C9���T�jE{��;�Cp�L��ԡ o��0]��$z�|����a����'��&ӹ���ۻ��_�����'��@Bj���&�	hs���'B`%�U��A�b`����f;�l!	Y��H���tS}=i�+!�h�K,��=��
L}ح{��E�+@w@Z� �	�M���2aE�Q(V�$cg���]#�`2Q Q���Gc�c�M�75j��������d�����H8�w���S9��T���׏�<f�2?zQ��q���B԰M_8%'�JCpb@�/���Zk��`�њj����9G�|#�R(h!G��9"�� 4��D_�=���k�K�Y�d(]�]O2i�N��"A���l���@�bR03��A�Cz��\9!�nǹ睝N�v����?�8�dx2�i[��3c��d�M�b���uJQ�k>ȕWG���V�3�as������H~hH#'���tbxh2�#dB�J��1�KB�T(zz�.�2�lB�r.Sп�������!�j���8��9�����H�6�#�`���[��~���S��;�v��g��bE��'J[�yBqÆ�Id�b��/�dg"�i ��نS�� �K{ȹ��t;���؆�;Ñ�������#��庫�y��x�z��xT�V�P,vt��S�&@D�����ly�UWm&EZ.A�sh�$�M�"�iu�ޫ���v�>�%�]\�hB0�{��9�B�͝��&D�,�ؿ�
A���Ϫ� _P��    IDAT�>.��&�'�<"P�L����Y�	������]�$�))^��LkV�T� �"�C�%:�*��H�T��=6�[bq���8�=�]��_��~� �T��;̪p^b�	�ŷ+�ŧ.=�zd�e��9	��.��L^`Kt��f鋴HbK���Q�8B�ԯH<�F��}���\�R�k�7���8A�q�a:69Ft8'�9L^C����.q�969��b��gs�1�M�ۂĶ@zok@l�+(BMQ�g5����R�C}y�-�������X��$c��)!]�S#�xT�0y����b)�~F5�r<6AH%_�� &��ݐ+��q\���m�z�i�"?v\D����� ƄƎ�=����G��/������O�/�~�3��/ |��3��169I::a�UIXlrv���2�$�?�|�:��d�:w<����O\S��	�z�+�p/I)�.�@6]˓" ��u���hd�~h����n��oI�K/l���ڿ������)�ԍ�L���a���߾��ǟx�~��[w�x�p��Bߑ�L
'�1[�Ӌ�Y��Bz�LN�-#���Yі�p@�EzE��+��П�@5fR��p�y]��PQ����4#n+��R�b��"�8xldӞvӳB�Kj�g)�&x�,UXV�-Q܏�Ԝ���Ғ�t�^����;u�:*xAw�J3yF��B�*x��j拴�gM;�z��������!cD�#�Qm�()�X��c��v wH$���Y&�5.���5�1*ؼ���u�L (�ɘ
DS��A�@�������^]"?�T����n<�:�x��
�L��h�L��6�m1�b9��`�������^��u�@(�D���[qVJ��-S��1-�R�hU����=7����α�.��:|t����-���������
҂�-�RZ�PJ�y�:EB���s��W����d����%�iʜ������=��CG^�F�^��=,�b>��!m�1�)l�~xv	Rº�w����on������7� ���4Y�b��Z�x��$X���QU8���<*���HV�>LXĲ�Iё�<^k(�$��S\�t���Q2�}�4<n��+>olU�4��" ��Pp�-]m$x�}���#����[\^���ށ�a�xJ�K�Ӫ��#YC��(zJ��Y8��ꕼ�S֜:av6�]hkdw���:�eg�\&eAG����L��(S�)�#�fLL��Fw��?EG!O4jVmP��pX���.H��F�V<��!n�x�r8�����6v���_8Ϥr�j��p�qc��/da��'�yFB�4��o���*�i�ob�Uv�9W�T��
b`<pd|4<V��4�ں:6_|�ʕ+/<�\L���LE�߶��'�:x�H1=5����%�V����G!���
ހp0�M�d��2	ev�L�_�m�#��4�u�p *J�r ?�	�{����i �%�kӌq|���nk�D�&
��Nl*Iǂz^2����i,�!�-�A��1n�Ǌ�f���{�!��C���(���!�$L$��B$:���\��f�PFP�uQ��d���?�ܻ�0O��rz2h��R=)�Zw[=	GzĦ A1f�ٞy晏}��s2�8� BR�(A�5[���d13E�(�$D'��`bۑ�=���d�,e�mk�,[��y憾����x�I7� �-M�/H�2�2�B����lF�p�핎v')C�:�Rx����������_�ȼb��J�<�:6ݘ:�` ^���?���D��Q'� Ƞ1�h᫟��0��3�r����
Y�y���SX$�f��Wɦk�v����prl��%� wǅ����Cm��D���2>��W�y��G��)`;\V��O@g���r����wHO�O$fӽVo�3_N[n���A8l��&|��%\5g3�������\ұ���_�����eK;�l@~ܚ�=7]�w�}�x��'I���'����/w�TPE�%�@��~��ы@�AB�H��,S6�y��P�Q�Y��\*{�#<��\Y�����}:�)v�:��ߎ,�s�:��vYWy��t��g�\ޖ��r�(�1�d
y�Ŕ�fs�9��:�w��h�x�������g�;V�01v��jt�� 𛡊��A�0�]��bW���6�X����M���PL��*�SL**ʙ�L>�P���>yER��(u�~�d��ڹg��v��gs��.�t���-ED��Gx�K�P��g:0D$o���ddr"�
;<���c�b�4)[�~��_��M=��rCR�*�aD����ȴ�Z�;w�>��K���O>v��N4��x�h���ɩ|+1�ǞAYb΁3��?QbkN%��U�]�ƽ��e�� �dC��LO�(����n<q2?OtR@u�W�^C�v�T7�i |��"�5%�)DL��S�|�b�2r"�T<<96T+�^�9g���w����߰�' ��'�t�%Æ}k�����{x�M�O�V�׹<��B��S�T֧�ҵ�r��\l�/]R�;�҃���L&b������z׻����t֦�0�3KNp�F u��.~�&P�/��7��o{��8z�Њ5��e�Ϡ^'�ؐ�A�A�	U�g�JFh!5$(���D���qT�4s�Z!�&��!�3;>15::N/�n[�h�'p�-���h�&������|����z�U�j�hxll�X,E��r�F���H��:��s�K�sp4�|<��5xl"6Yz��������=55�KA�� @����Y��V��{� 2�@���;c�:@O�:+DO�p�,u�8h5��sDV X!�m�l�c1��f��"��'p��j4T{���8�#�Q��ȗ1�~lt�)���hJ�419��n��L�HEr�=�A+,<\�'2��f������Q�;O芜����hY
��
��,�Al�>A�@���_}1+0p~�s��8������0��P����2ݹWO�wZ�*[�Qɤ�m�e�4�U�g�R�ɆuJa���G*��!t��_(��U����ћ?p�y���|���XoH�ogu����/:���>����}���p��o� �#�]�:d����xLR�_�|2�����O1;+%ɘ��+�I�&��N����9+y�jS؁��O�Ǐ����n�����_o64]|Lի �Vû���Z���-�O��{W�Z�˖ʲ��{�a"��WQ8&��P����O4I0�@FX p��R%BX�B͑-�<�n�0&����G�ۢ�!Z�T6�,��.�yo�����b��.Z��<�X�b/x�)k_wg��G�V6�qŦ&A�6�����K�|('IV��y J�Zb�/�� 24����db�B,��g�,N�Bd+��n���	����/�cf󀌺��	&DTlN�:v��h,c�,���J􈘥�'��T���Il^�`R`H�U)c�ML(���t��.���#���*��X�V�&�=�%����0Ca��JB�*s�B�\�N�ˉ+��"d�+�LnK����{�t'�c��5RYQ�'�T��Si��{!b Z�6�u��i-�Z*���s%�:ZH�|N����{�kyBO�˻~}��������u��	�f�7'������.i,�rG��h�.�-^*N^��k��7���4��U3w�V��e�V(Q_�����ט��o}��{�"�=�$���Z��ƉZ�M�}�`<���J�v��R���R����Z����ۊ)/d ƒ=]��X��< �ht�z��対�oY����OeT[G�u�΅�믿k��|�K�y���5�i�X:���˶�D�έc�;Ph���!aʕ8I�;F�U��#U.]�W|�DE�by��}�������@-��NMaC2�͛�dr�b��ALܹd>��X������;�S�o�@AN�=�H��j�X/޼�7_���~��{����>V�vQ�-zĀK�R�|`1���ܓF���#-_��#��Xsid=�7]uݭ��t�<zt�ᇶl��"���Iw���ѐ³���Zz`p��t-v�=K�����M�W\C� �$\?�����D�Hc�G��.���N����&.�TH3�9����F����%�gWe^"�����ר}��5&��N<r�X|cc��1��~��_��gV��a"���2��4��e���}�i��K�?��)�8�d�&Գ���,��e]�S
�d�,�)ȭӄ�^!�U�$	}1�A�I�Z%�o�喛;�d%0����L��i���Xg�����iˣO�'�!���Z�2(�A���WU����)(Ds=MW�"��B�N�3A��\#E�_�B�8�8&erS5b����@d�b�H��I�-�"�k֢�CqLN�R���8�q@�ΣF�C�W����'&E;nB6i *L.#'T��Gd�e�K�o����_������O��:<hN@ք%#��!���Iy�+-Q��Ax1io��J�z-��2�\�b����8�0l�ց^�(�5�dtI�u�MC���x2�
����ۭ���'Kd�$"�K��Nx����I�^�E�ב�U\�R��G�]�#DS46�.�>�����1��d������R�b�� st�sļƄD2��t��?���+7bY�����.ɦ�����/x���n$|�\r΍�zǶ�^�����'�}�L4�,N�?B+�C�4�K֥�qS���5�LV(1�h�5��G'FO[���_�B�{u�Gc&��:��6k��޼ȥ���f��׿�u���w|�S���X��4��!lB3e偲�"Jo*,{!������L��E�K��Ų����m� ��
Idն��-���@�L�)�M��pZgOw2���[�uǆL]�b2�tm�D���x�6�1����l��`9�[�	x+���[���*f�\=U�D��������ߟv�{^���/�d�O�ޘ��>�)�B
����V�6:�{ �f��v)P�à�\1�����n�����򽤵-O�FZ�ġ�ϟ�6E�
�Tܜ􃎋��f$��K;�����>��H�2bb ~e.
��K�J�)�[j5��Nʤ�S��4�*fA�/sR�p��ԓ�G�I�P7hQ����nipI���
���Zr��qth�\L������z�E��u,���8C�S�7��x��t�;H�}���O��*�Lx���PuMC���Х�����,ZP ��<ǎ�-�$�|*�^w��gt*4!��iw��iͬ�����R��=���&ҥ��'�\���\R��H����$��,���H�~���x���0�P�,E��b�nL��PE�R��b���.Z��ƶ�qX��+��,����p/EE� gm"��n�j��T�P$�<���7v�N�����l���������T6*9�6N��GR?�����Ik3�9�1T��������,L< �?�|L@xTUl'P�`���V��Ҷ}��D�]mm��A.nq���$-���튎���!�+�u���|�?�������ϔDQ��c�d6Y��G^Lp薍�����B�T1V�R�B������d����l�$�L���>���'�����e�DF��
]���;��z�W���� s
�8.�D�1[�鄠�?��7_y�f���DX�� fm���[XP~�7O��O��ޭ�m��/~#9�02Th��+�l�6LW�Х"�}��Lcy�;���$"$����������{��4�%fS�Y2I����޹�	N���|�J=��7����?0��/$h'[��^��k��9���O �z��$KO6�$ʙ�_�^t��^���H��T}~��/~�˗_v��o=r`���0���#3�=U#12,�]��է�c��߽����'�5l6K�d��P��׼�NP똣J�p� ߬U�����!�ǞI� ~������D�N,?jB���^�Qf���#�ua�\���md�X�D���.D]�6�Aj�����z�jl��m�����淾�"?��СC�>X�k)H�Z�	�m�i����H4l�%W�3�3M>�U��	���B`l"\�Xܾv�x�pQ?3�{xP,���35xfU�{|�%��S���3@�f�fR�����EQ9뜍�l>�J���*I0(�]E}o�(�w||t��^�|�Ⱋ/���{�c���Ǳ���x�)��Es�X�j��"�N��x=<�Zp���ȹ�	M�}Jj2���x��_����>��#)��.���(0u&K`�Ob{C~11�S�w�}���|�o�K�{������t ^Cf��O���!G�����9����\���ѩ�=zt��ͷo�)lH!�5�ۓ�٢�]�g���{i�5� �+���򦚷R�[���ɟ�,�Et3Y� %*��0I'�/�����v�ۏuwg'�qV��]ط7��e+�^H���<�%"��Or�H�lo.� 6�Dc�'n��p�f�$8�wG�Q"S�a��*]�x�Y�+��.��+�NMfv�E�c4��!�]&��D�o2jR�4$��`ו�D�T���� ��$�ۻ���!d!Ymm$W	����E�@e�\���k
D��[��9�ғ+W�}�������&$I]�:&��f����bJCZr���"\!�ʫ.;��s_xq<61NV?�a�qb�2�gף����.z�jM]��(���VK~21�y��^vQ2�J�k�5�+�H�+!o7+�\��Y�7���@�xH/�[r�-���G���6'i3p�t��B�0���۠Tg���o4CR����8hb�7�M��\�����=���b�O#a ~�� �Pv4���u�;x�U�1�!@p�݉T�����^�ކx���.O�)iud�%� &��4AI��2�%�P�/�◢�?�A���LV��tx=~�d��^�g�"����E ��,��yM}ǚ�:2�{!�aX	$�����?�F�I���i<���D. �ta�u�:,��py�#c�l�����?��t����U�p�
}�|�$)=����	u�Հ����~����� +�d�F��ؒ�ҥN�p;E8��ȧ,�iX}��n���k	,��ǓNL�7\�aݻozG[�<(�8�阉� ���,�l��ބ[�\�ho���̺uK���w:vw2�d��t�cިР��̮�:g�K�H ���R
E���[��:����\v����(�W�@��
Ñ}f�μ���DC�����i^}�/������q����xo8c��>Y)-�4�?���b$s���g��dxh�;�{�����e��|��]Sca����̒�">�@��M�J3ɂ�y<��H�L�T]8�Q�ذ~���L��Á�y����~���6�`��|�Ɨ�a�X��E���C��T�$j�;�]�;�&��V�XF��Q��@�@|r���lU�K�U�ȃ�P�&7�D�,v~���ۻ<5<m��(���WS�@'�i�ޏ�q9�A�,���wzLq[p5}����ԅt=�t����t{���n�_s��^��	b�J��Y��������@�h�]����U������+����5y�����nXD�b1�ֹۡ0j~?��"q=fq:�O�֘-kQ1�I�� b)�+>>xUD�?�o�s�l%@ъe˧����Lgg'������lwI85�'���ѐ�F��H'���+ɻ�g5�#�/H�U�5ӌ���s�T¥`�o���ۃ�`���*�q
���j��d}9�y�MW�OD��mp'�:y�ؾ}Xi�e}�Ug�]�?hmO�;�/(� ��'�OE0n��:!�lGe�,���I���U�ʪ����ʟ����r�zj��?:0p��9��n��	vN�W�T�G���`O�t�@6"^[�_��_���<rb�@܉���%�X��DAޫ�(  UIDATfB��u�^� 1n���.
�	ޢj�����eH?%C���l��z/T�~�>���J{���6�o�WG�C�4T�w��Z�x��
�D"�C��R�*��	��JY��"�?��7������)�� ����׷����!����J�Z:S�f;�mf�.3)!�8Uhެ���A�d�T��q�Bp��u&����Sk�Ѻ�ͯ��壼�$�Hg���e'Jc��b���2�)&��b�`���R=�0��O�P���D*��F�v�J/� 8�E~<J%~���: ;+L-T<�Saթ���@�A�+�"Og���r"[�]B�zC&k�D{^> -n�� � �(�]!�����QЕ�W'e����h�b�u��~��N��^���]9�3:��P��b$W���CHb�X�5O8A��E�\}5�e�G��R�v)��B��r��Be`sJ%(� �O
eW��D9]"Pw��'��2��(M��K���U@0��PA0�`(���!���+Yͪ��3i���,Ī��V<�L@`�Bl"?4�r(T�}��pjF��W�=]55�,i������s u�wV0r@�Z%L^,�}�0_v���B�ܦ��i3=�� D��f��!0#�4XRB�@��"&_�e��$��jp4�E^�S`Xj���߽����x{�D�Z��E�W��ئv��Ƙt��`]C��!q���4�>~a�F�bE}��DV�屛������K���vyH��Td
�� J}*����]�b�ф}��BY�T�
5�dg�S��N|�#5(t�+ �9ʼ�t���w��1���3��tiƕ���_���A�I���	;3G]�!���K)�p�9Gx�E��鲚�
Ъ&�ƋD�X�g��q���k�#�07�-N�MC�|[��g��l��kl×���x���` w`��:\�iD�ŔLa�'�Ik��o�y�q6�.�B�����U�xLv���x�P	���)C.344��Lǝ�
��?Ռ�نLj��o�(Y�Α���g�B��&�z��Qm�S��
��&@�Ta
�����pV�����a���5�p��\@�UX0�ݝ)��	�tNQ3�5p�^��b�riap$o���X���E�@O�B ouy��ږV+���Q��KxPᶥp�yH��bޮ�-��r�
�TG�V���/r�X#���O��+���S��Js	Zf�p�+�o��>����f�lݪ:��7T��2E�!�f7 sI��%J�Ю�10h��tW֯�A���#]IB�cbQPo���ƀ4i^�ݚ;�k�dou;�Q�� +�{7���լ�S=�g�~
��~�D��4�L=)[2���(�>���iUf�KM��Y�����p�����;c��B�s�Xcu�
�%FՂ�Xs��?��-?
�8qy��X�w�{j��k,���*j��'�fn��=W`jVɂ�}�(jYwvv����H2���h,�R>�M.���4��D,Ո���c$b $w�+��Db�N!�7,�<��~ qC�fCli13������*��TC�����)y02��G���E�3�/�h�	�.�I�Q���ɴ���ܽУ�E�'X�~ƩP�
��/ {uEa:yM�P�m�XDLLjQa�&ʆ�%5>�-5F�G�C��T�w�>*��qW��P%j;���� N�� T���@����_?`Լp��y����'�V2!��Q����A���N����%��L`�܁c���۩�	ޑ�ı���+����A�X��K�4F�	�.+b�?���r%���7�a�$��Jn�ĺe
5H+��L�t�<�=)��d����}�P?rP'6�CBn���NY�󕙗ʽ���-L �'�t�<n��>� k�h��@bQ$Å\䆒�PXTe�'�g-��D%8�r��9��tX�6I���WSv�lrT�A��0�BB�	�����Ŏ�"X��>��S��坼D�[���������T;�`˦�"��p��e�H8Q�:� ���ߎ�f�`��E�?z!j+�S�x��XW�%Eڃ�̾��~�=ĂE)&����BB*)�j�L��y�Ho<����� B+�ǉ7�s�f?|��[w^|�YӚ�z��3C�w8�����=��0�Z~���'''�^�L�z�D���&��Ȇ�+3�u�r�CF�+�Ɔ�9�ȦW�^M���ѡ�Z��d`˖-N���V/9������A~�7W-P�����v@K�C�N	8+�w� �	��J��f��|�2	O=�>a� ��9!zb��I��r���LD�H+L6��H1�q٩� L�D�Q�9.,25��i(y�)K�`��� �t,q�������kUk4��x]�����0�:��NDvR%���c��/�#�=�F-D�r??
�&eaG�/�G����S?^�`�������t�eW6.���H� /I��ޤf!�j"x��Q�� |`)6h�2S�&�딣��h�T���!�g��<�u,~�V!�����l�v�ޝ�~��[����߼ɪ���pM@�^�X�XmV��D��{�TB������/[���ͻr�r96-��:�}����T^h^��֏�����}���X�����l��Ԁ���h��F�n����o\w�a{ل��%�!KH�²W���HR���&��X2x����eN��������n��41kTv(ʡ��&qd��7�D��B�T��|�$���a��QA��!�H3]0�-{Dm��բ�sJ�y�/�t�Ey�t�)��O�B�+�ݏ�c>��㋢T9�����D%Q�,g���3F��f�rj��UOg"0�74�S�y�, �3U6��J<���G!\	�
�0|�vcU�<��|=f��NL�O|~�N^���JU/=jB�6�\�`��z`����N��#h	aĒ.�2w|��������#$QD�F�4\zx��0Boز)��]�"QJ��#� z��CkR63���W��Lr"Zk�3����]������{�&����0	%�j�I�	�4
������zCww7�v۶m0�/�x�R-t�vW
�����<��s�{ύ~����Sctr��g�`Hj*�c��� T��D�e����j�J��J�����~����A��c ������`Y��
��s�C�sE�#����h��W���j����	��V��������?���S����ϩ~�b�'�W��	�]�X�<(�̯�Ѝo{[g������{�h?�)����a0�\0v�׀�	ڱ����zܑh,uu�=:v�O~�|�qQqL���	\{�5�6mB{Γ�͎��3�_����Gs���x��}��XԹj�꾥+w��i��	:����s���_�"5m���6p)�a[(l)��DQ��,�b��tZ�Rv����|?<�������ا�M������S�%�	EcP�G��k�7_W�!J��8·�$�o�7�̖휯��}Y<?	��'��ٸX۩� ���$��3����@%[}�g��c�����{즑��+VA�v����VP��0�A*n�ҁ돕Ԅ��/ʻ��-?��}xQ�v���7c��K7_q���T*�kH��fP�h�򗿬O9b�I���f5�]����?\2:��v/��=t���݄ҊL�ٳ���֯w��xH������@�d�f���R!��0j����ٵ������l1�=���Q��/�DW��W#H��@�D�|�YG�e֕��XZ�����Ť^�-� ��κ����!|�u��9=�i��.^��!0?��:G���D��f2�YQG�m�t"~��A0�9g���ȑ����Q�e�b�#be�����6��������%����[}���Vn�Y}�B��z���ٕ+�@�
�6��Bz�i$G0g���E�#�����^t�E�^{�ϼ46��0>Qok�^�fM��ɉ�>��T>��[?��� �5�f�E�)"Ot%b�"�8쎟��;���۞}�@�l�/��!Lf�;#u����,��j�B���ڲ�w˛�H�Z���z��:�lt�m�_�ϿT��k�| ��j�|�Y���A��:���r6�A��pzq醑M�&���������|EHx�BI+�,�9�y�X�`mc7%쎝�����w���w�>���y��%֮]��oX���b��vA��X�0�3�%&P	;fT�Z�ۋr��CGʅ*&�$��ebb�R&a_��m����r{gO߲eE����i&�D�1��J����<�����<�o|g��'J����Q!��hj1(�]e�����U0憐�~��"i�qG�k��t�G��T�d�:jkȓ�Γ�ٓV�Ƀ��i�[{^{#��٣��^����Jv�j&ѝ�H��Bv玗v��ۻl)���B���P�p31wT�-�$�:)L{|����������b�G�ƴ����U�7���o��J�ۙ˦��	B�)�M[�	,�^�	�D�l�j��ܰ���ǻ�i��Q����=MO�'N+A��gȥ�n���\��[?���τ`-�26���q������������~@��l*�YF��d"v���Ca�,����i	�-�|R� ihU��;r�Ct�n��Gq�iU�|�9��'z�|������_��ꗷ�����U]����ڿx]C��`�Z��"�v�D#�����y���A�ːO����]���~a�ʕ>)bĄ+B��`03:�ٽ����|�@,D��3�~ƙgTJ�}��R����D\�`�Z*#�$���+.B��Xa���y3�p%�ց��m��#��X�����F�����<�0����`�m`���]���R����ɉ�;�q�Ҟn�?].�aw�Џ��yj��?[,XX�=��enw����T
�H��G6��=!ޑ�[���V�\!T�1s�2������W��"�����5�J�'p~\��%p��h�|�:��	�G����s��X��,\}�LR�r�J�X�-��wvt�/^���ccGGA�%�#�~j`��|��V���N��8�S�b��wo��忂 �@�ښ�ַby$<f0/��/���	���vl�*����+U�%�*
�4��	�	�x��_�z���^�P��@��������fK�"�Ap,q~KFbVb������	]��p�}� A.P�H8p"��.q��%1�l�p�ly�<�-��BMj��a�N�lh����[�g�����[ÿ�D]|�"� @$���r�Q18�G��	��ų�\&C Hu؆�� eW�P�Â���)�=]��rn|�h���V�[O|�/�>U�$^��T�ꠓ54P��	��.�u����}?���綃��%���T<�s؉���e�����:�(cP��!zI<kUR�bs���C�M�}�*�w�H���Y�=�>�c�N�)��Q�]�)9���oUN���jY����P!Ц@\�w�:\��P¹9юH�YBǦ
:rb�h�b<$~՘��]n��.y���Ԏ][/�x��?���������ܬ���$5�	Ҡp�"�43N�hRT�6Te+V.�hC8>�:�T4f�a#a�m��0�m7:�!�٣B^w��GK��O�V	��wy
�JEV�P=q�m&�:���bL�܊�s��o3'�ʪd��k��>�G��4���o���X��+A`��[��U*И,�ºB^0�rXg�Z��0Y�Q��6����>q�ݩX��5�X�^3z�����/P�B��T�@�%f�V����?̃.u��t:��3Oo۶}ph4I��u8��$�9$���&W�+���E,6h+,.��$�y��G.�pK���ICD����ĺ�TZ��F��{7�䅧���jY�|����ŋ�X�@Kh|���qQ�2�fK�
�<���$u�����?�j���B�R-���`ghÆӗ�Xr��uW^��3֟&v�}ָ��6M]��"65QcٹH3WL�V����خ|���x<:���a����Bn\�n�b%��%�%-j1�%2��9���4�u�UDl�ͤq@|	�|JKsOŋ�cU����\���ih��q 0%�����錔�\(�Є���&�=F�Z̏Џ�m.��5�&S��}�[��jt�\+Nu'�&�',<E�C-ī__�9�����C�r�fA��uМiblrﾗ!�K����Q�x�Pʗ%ܕL3�#���A���z���#=�*~�Eq��qc�u��U��Ve~jN��:٥xP�*�Qǭ�]�����o�J ؆zG�)��A^�k5�$��o�"��n&��P� P~��R�d}�Ҟ��$%�Ц37�Ͳ�<�B:t�TR�.g�K5.�&�l�X5��务��R&ޫ�|u�Ŧx	�*�2��Ġ�&F��C�����hD�VI���P3+�j ���!��E��j)��`:�f�#��@�I&�$�
�>�b�(9�ȳc�J>r9p�A�s��Wt9ݎ�z�;3��	�QǕTG�x6���B�4�BŖE�M>nb�	9���I�][�P���R.�z+B�R�bY��"!0/��)�*�.��ʭR!�^�"d��@T$��*6G�29V�9ېI�w�4��\9畠�E��8�,^X��"!�����K�X��"!0�Et9�ųE,B`� �Et�
�Y�i�X����,�!��E��?)H��=�O6    IEND�B`�PK   �x�V��K� 	� /   images/cd1eebff-8d4c-4172-8358-6f93b12ef793.png V@���PNG

   IHDR  }  �   ���    IDATx��ߏ$�u&��s̬���_"��hDZn��� �o۲��4���/k���a�w~�_�I�a�G?�����&�ZY��"���RI\��a�L�Ȫʌ������U]]���=�3��}+3�Fܸy���q	l��l�����k�?,N;�|��8�l����R�:}쾺w���=Q��O�A+�{�p��ݍ������W�컗o���4�A���Ʊ66VE	3�3�1 ��L���|bwG�� ����E�Mk��`�c�T�fK�<k;���. ��p�<!�ݱ~3M��5�����6 $�� �Il-1��h4�a7��.��$��)�ԕ $����9A�:0� ���Ա�x�֭��#ߍ6X���`�VA�e\�v:���W��l����O��TCn��>�2r�������yf�/�i绺�G7n�:pف7�x��4�8����W��*� p㪝<���ת[��������1p]q�j��]����󋴽���X^G�S�G]�X�}wkw�
9�nW��n�k�/ �_�s��?����l��2� |0����h~{��v�Wf_��ӿtܸj��օ�D��Cuk���a�l�����f\���X�{�u��?�[;��/L;���_����z5`�Ez�ƴh���K�H'wk�����bq� �`w¹=��k���=%M-����|��&�k׭#b�iD `㎪v� x4�̈��e]s"	�睙���6hѨb֜Ț�4' m���d�*�Â�ĬaȊ(pqA�HJ*Mt�5���B�f��^�֑��X�Ξ�� �)�8�bĉ��OeѶ����,���[7o���y6���!}l��5��=�ғ�a�m�}���)��bw������-(�)]�-�i�`5O��#	�[�)�w R{��;"4<� �6Y�������wp/D ��˽�ד�t��v�Ȓ�R� f��(��Y\�JnJ�.@�EʒR�q��C �� �$Χ��� ���vN��Q2�7L�0ClG6�����	�g��{��>_Mp�s���1kZ����m�J��I���%�� P�HM�XP��5�&��BV�e���u�6k8f�ց_�T�u6��*�͕@]��
��4Kpk2@L�LFU��Ɠ����Z�"8 t�� ��YNۉ���'GSG�G�=O4����f��� ���i&sj<�mQ�q�g"��a�� i!\+tЃ��`�Ľ�`����j�W�ա�\ p6�yE(*1��2���0	@Y�j�q��gU<;H��nr �܌HX��p
�.��s���$vD�E���;XjZ���L��Kp�2A��T�X$����@�DN�Ⱦ �]u�ZR��f֌����o/��ݽ���p����|�!}l�cUm:������y�"���M�tA�BKVg �v��dm�Q�	 (Ufi�j$k��y���q�j�$!x�����.$�<�@��N��I�R�Y���C�:��Db����8J�kEu��"ޒ�*�N
��)~��-u0��F�+}. ��%q#� A
 -w�<">`UE�zb�j0��J �K�	�]�,��m� 0� ���8����$1֛�L#�*y)��Lr
�6��+ `/����� �������o3g*���K��4j���fdB,p1#6@�0Aۗ�3y&
�uq3�A������ȉ��!3w�35�fX�laf�1�HJ�89( D�D,�Np0*7�	�
^8�1S�1�_��Զ`6��#0܍�����O;�����[�Z(�`"8;� b��#r L��;�`�`q5��s7V�����sbe��`'r�	�N쀁�H]�D��0�3�3��RZ�؅@D�09��	�n��@p����F7��0� ܏���Cs��2��R7���_Q������_�o�����gkU�6xHlH��k�P������u\[�e�n ��#��l6��t��z��~�����eH���l|)H��/��t���\�[��Vs�q��W��v߸���׿Y���y��W�~�P����E1{e6��f^U��������鬻��� ���Oo������ʕo����On�� ���6�{�h�s�;�=':�;0 i�"�Q�u��ig�Uv�ˣ<ˉC�jO��խ�LRp���dZ��!�LZn�"�V)զd1RmYTr�,�� b䦤��X3s��������,,Ɉ �F�E�č��؜� 5�T�M��Ɉ؉p7B�.�Q`!� pa 7�Hԩ� R����ȸa�ƍ����Bd��I 8ca�#n��HU�*�km��NRiCw(��``("mXi˴���fi�Nn��d�7�12KHn�q<y[�@��n�R�9�<.�.�Z���ͣ�	1س�XXA�P��!����ȁTc�P@ b1��"Av�����Y�FB!!�`���6S7 �X21��3`�&8���� �r�@@V%*���ЇBDH�F �b�;�PJ��>��/ڗ��9/��{� ��X���D������%]~��%���BVEd9��&�����Y�DC@D`n���B������!�CX��>�Q����]��n�q@���~��27�aC��U\�����/�'��ݳ�싴XܦU_���6��>���C�����Rj�mƥb� �[e��>���{����lF7o~K�\�'r�������7?� ��Po �}���-��Ɏ5{����3�9�:z߫��l?���7��x�Σm ���6 pIw����kw�_�A�\�Ej_ݧ����+W~"7_�m�߄��7��ۣ���������ݶ�"\
5�٪�ȉ�N�|���G�Ż���&�CUo�t2��UK<χbR�w�I�B��#
 �/Q��(��S�J;��[ud ����/0Y�^Ea ��H͹jY�MI` �$�Y���)1��D�b�\A��8���ڲ����K��Y���q���q��Dn��T	lDfS׼��;3�AA� 2搌� �n@�n�pb���s�ى�����48,�A�M܉��9iMd�
n��V�1p�C�e^'"q��9P��R?/ܼb��j$��H8�~:P���{����rm� ة�O�;ء�B�@M���RO&�0d�I�	 ���ݝ�(lD���{S�9 �Q육؁�2�A��L`�
��s ��[���v���,�O�L0U���
���0@������(�
f'߫����0QO��i#��`�c� 1AXp8?@�����f�5"Z!�=��^i#�e�$h��| g�*��,�\U%x6dS1BX`pXV�	n��@� f�!<��렙A!�0xT��9�Ӻ��o�U���|�'����_�c�΁�&黶�\�t/��~�3����+s���6�?���72��?`�8ׯ��.��w��]��b ��4dO�J�/K�����ɓ�ҜbyJs��?��v�"K����2����fʾȦ�8�X��b䣼4���#�"�(Q�"S�r���X�`ɫ�7�,�w�u�h��� 8|���H���F�)%WH�!���� RU�P	{  TIn�¹�N# 	QɅrE*�kVQ3M̤s�A�j��HsD��IC4�6xb�3�A}T�`�fO"�N����F�n�U�p��斃��H&h0��;
��<G$���5;�23�č�7
�ɼ��kU��y��F������*3،YrΩ0��0��E@+&�Vۆ��ɂ	�ĴTZ��32wv�ѲW�]t'&עx��̉�b`w��C`�p&���d)	4�D�j�n8�9l�T&[e7���D��=��%'XN� ��hRf�^eY%Ǟ��{wGUU+�Q?�ے�/�wDhL ��u-��	 �p����#�yIrt*!q7XߦJx�"���T�( Y�����/$�
�1���?�c�"�9
YY�VK8�xpi�ɶT�B���)d�Q�-U�Ổ3��~�����BX���!猜�{Z�VT9���ѳ�~��po�^U��OwG��^�#�  �䅺y�_T��(��̑�r6�	B�Q!%�dk��f����u��W��s�YS��Y�3��[/6��Q��"}W���G#y�g?3ܼ�_��߿0r�w&�%�z�/���^����o{G��cכS�>�jJ�> LsG6I�yD�q"��J�} [  _tc�0w9�\']��9B�DHt�ف{�.k8O
�#�$�$�����] �ٲ���M�?� Ě�ݕ܌:�	�z�P�t�v1�aQL{F�ܤ��~���9S�W0�\U�8qq���. ��� n��+7ew'rnĮV;�ʈ�027�I�9� ��X��lv��~���f^���5��D���>H�>r/�WNNH�N`�5n֐#j�v���LD�w*�+rSm�Zkֱ�n��&���	d�bV-�h��Z/3���݋�X�HD�� D]���̹�W�݃����:w��9�����Lp��^�A�A���;�ɉظ /Vբi�kp�`���(ʒ�����'DH)���w�O��-KϚY�T{�a��B�{Ť`��7L�,+�:V@1��RiԠ�W��������3��$>"Z'�Ĳ�I\�X,���DTHM��b�0� �ݠ�@�7K�k DG߇nI�j�@D� �z̡��H!J�<'�d�)�Ua�����~�	q_�=�	N�����B���Z���C�ê9���K̣+fU@���'kǮG�1�x���`.���'���\�4f�۶(��yE��e�����N{I�<�������c���!Z�3\��3/`�U����b�:�(�Q���X�3���;��z&vx8�=�y�鄾w���<�l�A�O�#\�*����y ���$�b
 l1r�NA��F��Rm�L3yUQ��r�1��R��*5J�Q��:��SͰ�������H0{K\���8�{�F�L[IiˍX	yf��2���p##�A<� V��=O�hDN� �-�_��TGL��Da���;^�=3sΑ,o�c�=m�9���0� �+Sq'*N?%�s"	3�q6��W�:�[e�FnV�Y�Z݈X�qK���qf�� �������� g�VnV�i�����;@�O��DJLF��ff�e���4�p h����Ǡ�Tw6w�AV w_y�/e�����߯�R(�G���į�8jc��o�-��1FQ/jUOO�W�K:�
+��)P��#�  ���K��o�R�)�$a���$���8���ă԰�yL|��	���j�Q���ĝ~��k>�7VIV*��Cv:ξ�b�\=��,GJN_�J���Y�����R~��{�p?�z���'{�Ҥ=��} ��'="q'�8p��=���B9(���A�z;)=P�$����7O�8�p��u�]�����<����POƷ�i�|��v)��໢~7v#����?>W6�L�&}/~�7'�}�ߚ_��[�ίx��&u�'��nF#v4��0	��]�Φ���6f0�=��� 8��8$Np"U�"�)�m1s���%&f%|�@���u��P�fp�LN�`��Y��j}�J Nŗ�j��Ld)�F�1���C ����t0�N���U@�wJ�ٜ�H�wg7��������{/�2���SQ���c�Y�Y��ưB��Fn&�ΰ��Dȣ��+R?S���/�Xg��8��RQ�nK����v�� C�W�C�ɒ�D�_�ލ݀�����,e��� �z̄�z��������V
�Mv�o0	�lP3�X��٬�f>V���=���|�oR�9H�?^��ޠ�4v�p�$�H�2i�������K��c�ԣ���,�dk��_O�ζ���okHǺ�����{$0N'C[���ܩ�ޞ����>K���pd�]U������I?Y*���[8����pc8�5�F`éF�lc�X@I�!̺�EB���p�;c�� �8���[����o��)N�^�����jvv��o'��v8��g��1"�L���Cĩ۟o33�#S!x2*
���($�̂�I�/����
+��Ɉ( 'b#"��<�*͹���dfK���`��o�ۑBS���(RE��?���BÛ��3p.��y;��2�����j11X�L_�ļ<^�BsK	q���������K?U]�9�<�99�嚭?����Z��В��1I�8YS\����f2�Q1��Tw��k>S�2�/���p������P[�A#�\W��-o31�m_�>N�xP��I��0H��'f����VHn)Kލ�H�~ߓ״����u��	F<��~l��G��u���={�ZR��|vm@��i?�|���jWʓ�����Ǖ�ӈߙ��`���-�bZ?��wZ�����~;��BO�N)A	�!}�ZL����@4�*R�Xd�֣�k&�;K[/c{��!ϧʹ��ǿ����`m�m��a��ʕ+�W^�V���7*������~��`ވD mآ��lPYV��l��T[��ӑ��ia+�F�<$ ĸ$; V�8��t��V�&mf0�š��b��Ӿ'Ho#�S���IA. {o�Q��۝A'�*F��t">Rݖ�G�h���ݱS5`+oĞ�e �� ��0�2�9JTa��&ͶT�Ыi0�3 ��5��2�r/��i���i���v���
�^�0�ș��i
��Q�{�nu���W�_U��O�A�r�A������]�OW0_�n=Ni+�`�S2F�����x<�w������jI>9��k��s�YVR�<�yW=߷ߐb夯�i��)\�|Y���*J�����5J�Z���g]I�v�ώ�[�BBP�U��z�������Pwp3�����nF��ۉ�;�lr'�r��o����T6���T�^���t��֔��M�e����<G$�N��en��];C�4ݛ����+����+���g���:�)��8d�8�J	�2����8�s�����L, J�'�P��86�y?Xi�X��i�{�� �B��p�\��J�C��T�ݏ�5+��I_0 �37���6�,� (�w�lH�� �^a��|٧�  ʺt�&/�E�bf,zG����������~�tr���}߭:���!���'�=Y�>��`�Y-��C}*<���SQǎ���)���>?p����q-�u���>P�}�`�U��)��ʳ=��W�>j���B��o�����K�?�D����K^s~[�~ZS=��~@Ik�����71� ���e"��>�al���5Gj����9��(&{��F}��z�0Q4a�?G�b���b,:C��j���4�݄�37:fN�9�����t�
�9����߬_~�VuYh�}=x���E��!��!'CUai"*?|�#�����:KW|� (iQ,��x9^*C�������'/D0:!�����	� �!��2R��p_M����&gD�BV�$w)`}`�����܏���g�c��<~�t_�-���A�S��>q�w@� !�rF)iO�2  �s�{��4���<곤�Ẳ~���~G�vX�!��r2R@��>`���_�{N���QV�J"Z:嗈����X�����'�>��+���K�Ø���K�����$��9
�!��U\����W�e����8�(]k���9?�R���!�]��T�p�Rut���]�m^4�3��5�זkH咉= ���e�=Z�b���!N+�V��P꾟���r����~8�qQ���\y�`���
bU^|�6P�Te2�q����<n��ξ%�e��կ~o�{��]|��L<�x�̻����zwwk2鴍i˃��5����v0kǮ���y��C�Y�E(�Tn���1�ʭ�C�QCZ�..��X9oO�ZH�z.����|eK�B%����0Z��R�A�q����=v����Y�|r{�vi�<P@~���~?�C:�#��Z���)���{U];F�؏)pG�6x�o5�jJ �|�OӀ��o�߸f\!���������    IDAT�$��8�ϱ��ȼt���z����OS?W�'�z�����'�,��`�����a�~������B�\���lҴ��2K��Wa�H�٥�{<�E�.	��~���#z�=�����pߠ�Rڠ�?h;1���e�%Vp��� F@]�`N0� �1�@�����i��P�I�OM�Z������}n����ި~��3D���_���Nr;��h��^|���^�����k�qp��)c2ق�G���Ї�a�~q��Ѥ�:��䬧�� "䜗~|Gj-#�Vsku���;$��$�p�ĺ:���l5��0۲ݫy����$m'ɓ∤�cqL?-I��>,1���պ��|�uߵ���6�"�Q*N>�m���A�?|�S����m�R�c�5s���g��a��q닝��܁O���엎���|��%�{��u)O�<�8 ��9�C���}���x����֚�g?߶������� 60)�2� ����Pw�W�8��$0`��jBA�'u�C!����p0N���}p��� �!���o��k�(.���H�9����`q�+�Ҵm�'?EY�F"��{�=�p�nE�s��9c�"N
�`\J��}���&���������3��úIeݠ�I�yI�:���y���4Y�'�,>_]��u���دo���?����>z��mI�J�w�X�Dq{ƶ�?���K�i��*!Lq��tuK�?�P����0S��������n��o���ݟ�4��;� G�*���V_W_ކr1�0�DwS=��t��s����"��"h��߿{�֭�ǗO��3Y���ŗ�~���/�Qg��������TY��;Mڶ��8��3�w)Y�w?=���P	'�/M@�O��q��� �Xg"|�����>}R����<�5}��w���d?|�׷w�NN?~�Ԙ�(Ռ>�h��j�<<�'"!,-UU��k4M���QU1�Ǆ&61��
"		���7PI��N}��@(�KAd�H s!��~-�չ�� ������j���֎����*�q�ɖ������9���Έ���_Lo���F�����ة�EWј+{9R�1����·�;<��B�G� "ǖ@Zg�|�<c�ͭ��཯��D�2��F��A�^�}>��Ügu0y�y�{<;��Gy������q���8����X�2Ƈ���@eUA����������R��ޑoq��_�w<۝��
�s+I�ѡ��g���fF�]V���SXv$�% �J �$j��Q�FK׉�����Wz���3>�ן��HmB���l��E
���D��.��ю���9�7[\��\�ݴI���F�._���4[)3�_a���<����T�"�Ï[��V[��*���`K����zp�J�;�ez�#��u)�����I�����bR��O���?��u�����V����������ó�<:
�)k�:�O�>X|Č�nB@UU��
�
&,�8	;��KB}%"\�
�sԁʋ�;̙ �LMܝ��9�,-/s�dG�Nd�rMc��7��c���sAoI꯯���}��yI|sF���6��yֹucS��"�#�c�x�vƷ�`��	��,�'}׮	�_���[ �mH�F��ۃ�����ѭ�؇uC��R�;���;(��2������qz�+eyC%�r�9K�{R��*�|p2��4���a�ϯ��X!|�#ĒŬ�i!5��k���T�-H�8�D�2�1�q�T���"sr'"cH�E���%_1�G0�Y͂U���!��S]J<d'�`���,�D�S�/h�XFk��y�L���� kA!T�b*]�9������,�����`�{/�7���?X�U|�O5>R��+W��Wn�F����	o��z�s;��������l7�L�@���f�$|�
�O��9ͻ}:�eb���b��WV�~�C��*���M�q��I������I7�=m|܁�h�Q߯���x@�>�����r�֑�cfNT�B���	������������q����B�ma!̉E2�nj�Djf�UM-#e����]ۉjY�@�ܞL�D�����*檪�X���bfFo����^�t`u�l)���ݾ�Mj|>�g�,��U%x��@nI+&e��]���i-�+_����5k n�i�GD����_U����2���T[����?�n�w�޾��f��2X#�t�-|x�'a�%�F�jC�MF���� ��{q����sr����r�=��p���"~��?N��iWK���}�����G9�3��w��������n����W����Fy�>���c�d�`:ckk�QS�:ƅHh�� �j�9+���������fN9!���Y6�dj9gqgu3/Q�啟lC�Pa�����2sF���AU�,B�N}ri���,��,=]V"��Ւ?\��m����zOЬU�d�� u�!�6g��Q����^y�[���ؘy?�x���+W����V��ua2B�������t���������9	�W�_>��sFJ	A�N��t,��1��P��J2cC?8�01�oOg�|���'}ܳ�I�78����5|^X>
�>��ݫ}Gc�t�U"oG���4�$	�� �W735SS�;����)�T3g$r,�mx� c"���%rd��ȍ9���� �  �3S`��Zq��@U��s�4U誶3tI�@�'�a(�C�ə�劉}�V��� ��VҘe#�T�����dg���>4���D�ݽ[��gOqd�&_��_��\�_���1�zȵՠ��ٝ������c��R:��w0�����
�y/��.'8;�* \��J0����|�n��r.�idYY�#3��Z�+H�ݔ�PZλ}��yq5��<i'`}����~;���i�_���i���y�i�uJ��Nj�۾u.�O2�H�^R�ر��"��7l�jL&4�������%p���	��[#fN #��	� _U�7�5= ���vx+ �|DBu�p�1��Y����تCU[j_��4� �Ч���*
��qN9�9�)�kS<�/0o3�ڤ��� 3LE�vƎR�6f�ˎP��XCUP��Cr��A�x8j�w.=�'Jp%��o6�_6��N�C`o~������3��������"vQI�y�/՘����蕶;����V{0����)��� ���fĩC�������u�瞿�K�.a:�b6�������w�.�Z����~zr���,89��~^]x���6���bu��~�U���fAU���5B]�V71��SA�ٲiVPb�d$���C�]��D��s�w��]�n�����s�������� �v�����?���k�x�G�ɔȦ��9���5@� "����R6�='!"&�:�ZוrS��Lc'�!d��?9 �e�P��8�7�, ��5L�բ�	b�ȠI�"�L�*3`���܅�����)<i��_�����6�9F��ط���]��^�ŝ�Xg��1?����K��]Y�k�,=���Tu�[Q���f���~�~/�������������],�8Β4:֮U�)y4���rR���n��''�#�{i3- ,�QSa<��:��d���]���)�Y��V�_w)�����_(�w�!����Y��?���iFYj���Kӗ���3��a�ۉ~�7S�������}��H��=m�N��*[�:����/��9���McbrS07ĸ��dA���-;)H��'�]�$V�;�Go�-���(��()窊�0������bz݉G��ҿ:����'I��K_�&u�c;a1�)�4�2��^�D/���7ݻ��.u]/#tO��V�݃�y��䏙��(I�U=ťK���W�u���..=?��d
!�Çڡ]d�ԏ��A�;��s� ��i��6�pޜ�R9!@�4>]�=�ow��g>z�x֯o���#j�'O��a�op��� *)�����4�WU�	�"��H��J�� 㞃�5���?���)�Jh��q���X/|��<�ߞ�m��u���g:�N�ƍ�����ڵk����T���!u8�����O��>�į0���>�S�m�6����B�,�w&�ö����:�_hZ	�x�~_�	�}(L�M�$��PW�Uu%�źr�W]����ՐfѶ�	��≑�˗/ǪJ�h�O����\�ؾ���Wg�����/�j#��k�e Ūo��7�i�w	N@
�x�X&P�����jR��C�w�{��-��a� [��4����ն~�m>9	��g�7,�4�PUT̌�|��_�w�>�89�G�_y�+/s��59��s"����:'�@|/�����2�7�����\U�J����W! \U6��Ӆ� pJ[���<���oܸ�� �7�x�oݺE�/_�7�dŽ�_�v́��ۋ�sU�D���������_��k��M^��?�.χ�_c�_�L}������Ȗ���XJ2?,��@��F�����S�V�gAq�����8U�(ֱ�+a���+�w�t�]0���+���� �T�z�ˣ�횦��4����(��������ˇ��/T�
A"rJМ� �Ӄ4��qe�|�f�%|�N�!�1�z���Ӌ�nM����* �	)`1���|��v=�u ��x$��9�V��y�� ���OK�1(|��[[[����|9�e�σ��qj|܁Ow �:�W�{ځROkۿ���x�OWD"��H0OP�U�U�@�ݡ����3�����ڬ`����������ٍ~��^��R]�	���,�(�5��trX����4�F|�+_�����o����bs����{W._�������ƍ �/_0q]���_��=UM/���sq�"�����O�v5���:�QMG]ʵ�s���3sf"g@f
�$>��a �%�,$%P��!"�5ƓI[ג��S�uf�����J4����������-�%<�w�ʕ�4V��Ӧ��RK���-�����K9�q]���03��s03�FJ���3�z�7�)A���8ߠ˜a� � j"�"�d%<w�yT�B�D����A8!�C���T;ޣ���?���u���?����^�F�P���mۢm��ҏ*��Ӟ�?��i�_���9�����������=����5r���*�'%8+1w!63�|Й�:�/�eN򝪵?�������/��k4�ϫ�~������b�@�Q�9���Q��㺙T�d�ĉ��gf���Z4�{��s�����ޞ���/_��/��������������/��a�ʡ5�f�R7�@{ �CgPG����+�Bdf��vPSD$
��㣌�Ď�$]@VI ��q��*����HB ��kSp�Y��W^��t6��͛77��3�'B�&�I|^���V]�"��|v��pߩ뚘�Ѷ-��1��l6�0�L��\q��Wp^ҧp' �5�"����h�!����q�x$ :�3��[3��6<K���i���>�n5��d4���z����������=���=�'�t<����񒾓/t@I�B@�IH�,1	s���~� ���?0�n��>�����ʅш�����l63`��u-�k"��@3��0�ɸ�Z�!��
&NW"�$�:�h�9�d2�w�y��|�M�|�2-�L&��/����� �����o;���޾���Q]��� �Ax?V��l�97�5V�� b ��\-2-鼺sN�D� p��8�����V7�k���J�����[��ao{���×�Z,���9>cx��~��~����1}>��_U�WB75-�/�/��@�BN����7y�,9�;�fo�%��̬\j�D���dG��Ü�0#s ��SꯘO�r���#S�&��!d�[�=+��×�����y�gT�R�,�����#��m��}���jl�ꉦ�K���&�1W�8�ZTŐ�\~Y��Q)PM�u S]{����,"n����2&V#��6�r�%��.��]&�]��QTJ�Ή)PWC����nd$��"��su�6xR��c]���\93#Ɯ��,K�?[�EO�Yz�΅�w1I,Hߢ�岥�v;�:~�+�q�h����<Q~M���Y*ۋ^��B=��̞�}�=���X�w%
�v�����%�v�ųr�˞�����Ҿ����{��O>��%;��by {�����%���E�i�?��?��@K�����-O�QR���H��tx/�W+�+U¨+�ՙ��KE
���_�ݏ�[���t<�:쿴9���ɿ���_������+>��Ѝ|c�@k���S�2UfV�5X4$E!�h`S@C���A�3���,�=��g�{�=��?�g<x�@���x��!�o��?�) K �ө��_���W�������<)�� �w�ӥBLDER�O*t��#!�H�ǻ@̵{�#	o���pf�D�%,u�)\IJ
�����(���r6D��HrZݼ��&�ϤM?�X?��%����X����˕�~8�x���E廱�7ۮ'�.��B& �W���D��D����50-)�cN%S
��_@����ӆ�٬!�D2!%#�\�1Gg	}1ƥ������:�����UbA��[��[rGRۉ�}M��u���ܟ�F�ğu�g���'������/�ٺ�P?�{�>DdA#�iۯ/�^�1��<}�_�<��~��Χ)�2��倫�TQ���pYԃ*y�A(�>�r�D�؝t������D}X9;�"���r��Ϳiy/w��`௪��"U��R����
s��`f1�yT���ټ��ҹ��UA]��VA��Q5gÿ���2���{v��m>���Nj�ш۷o��۷�ʕ+:��h4���?o��"�,����R�w���'j&�L��BũvmG�h/���q��0lH_��l���)$�/�IA�W�F�4ճA]I=(�:_t��d�KH���\�t4��}��¢w0�Bw�B��l`!�E��2x�y���G~�H�耖���!-R��z�2R3���|�5�7�"ZҴ�vi��ug$b<w��J}s�Χ�Yv� �d�_��"Wy��4MKJ��)�|��_�Ó��Y��I�+/���� �.|��=ksu]RxD�s޷��M����[���ck?�+{����z$�f�SR������ӔJBU�eт�"&�m��Sl�R�M:��������������ߗ�÷������EU)�g�B�`�y�y�=tg�}=9�& ��]�����דɤ�'':�yY��ʪtq�EIm���w�N܉+$,qJ�̈́�KOȨbNI_|�RL��������*� �lg�}���}�/�B���:��0��"�(�T`H��,&qy���f�	y��b���8j�D��'�����{w?e0t�*��`c{D]�ܸ�&�yG�%��I��LL�I$�qX&{�Ƚ�ҩ����fvj�[�vAϓ�K\��F�k�?�\�������W������8_cvA�ʲ�����w"�9W�!Y0ѓ$|<����%~��do8�ι�?��4��I�O.�$e�K�Ue�4�YJqn1��Kݏ�ſ,����4����O�@x�w�w���n������M&p��������4�`�B��/��q��b[&�J��ŅXk3���tFJm��U�ˀ�����L=�o���}�YP�d���P%�����v�Νˇ��B���@uh�%+���>S��0�I�R�\����_�{WLs�Lb���`�i���wLg�|����XU��
W����u�̛�d�2o~�����
e1rZxmlp: �w��y�ނ�-��2��]`Q��-�2������l8��л�W�����$K��ئ��EMQID;�4$$$�6L�毛��/���;W�p6Ҵ2��h�r�i ݊�t��u�d��*T]���.���nA������� ����ߓ��=K>��]93��F�k�ʂ(�֩�#1)}�����fBe!�Z����D/�-�������ԏ���	d��B��묒��=    IDATj
�����%~o�"H�Tf� �@x���8������'��'w�G\~}/�mrܽh�E eل����!%v�fT�x���Y_��S�V
VV7�q3qp8�`�������]��Uw�#��	~� ,�<_t/[/.�Ó��M�|ON�l���}A���,}����x�{����eq߽�e��"��!."�d�����>�7�_:;�����:�IUuiY�~�e���(��Ƶ����n��E�я`��+{�'L���hu�b���9��]<��M�Mև�+���z=F��;�R]U�h4�)��e�Y��S�ŔT�,�ixt�\�Ϟ[13�>h�""`q^J<��[���x1�]�:D�h�>�-O��,}O�$�����D�.�jUI6�R
�����1�W���HUU�llq�֫<x𐽃�>RՈ]`y@�&R��ћ���� �ǉ������$8�:�����*�|����-}$�����,Q�9)�Fq>����ʹ���tP��u-�9��,'[U��%1��AV'���7:޹����v�������;X-�0����ae��}_���Ͻğ�����m�d+��j6�B5/g�]ȁݽw�=v�x��]H����0��RBP3K*�daݻ|��x��'`s睈8�d�X�3�>�����$!�"��\GY@�L�{��~�)��̍y����u��+����d82�#�M{�."|˯ǥ'9M)���ey�����%~��h.�b�u=�^3�)����R��y�m��]���ڞ����i~ûr�T���Ih���������	�N]�-��Ģ(���l��?���pؑ>��7�~��"�9�J�5x'V�SAI�"��;���v^���B���B����bT�G_I�\��/$e˛7w*_��\�uD^�m�>�M�'�$�47���I��`�9Y�x�;pa2?M9!��֧QE���"�*9�`��%���
�j�`8,&�M3crrL�-�tc])\AQ��m����nҋ�$����h/��-o�eqQ�/���c.�^��E�]��,iXvO^�%|Z_[>��sXN*������'eٲs�<����{s���y�e�ڦ_7����Г��Y������N�~�۩#�<���+��K�Խ����}R�vP��	�!bw$���l��]4x'�t큨�aR
W���b{o8l���w�?�����-�?��]�r%m\ۈι���w��^��~P��4�:�𾬮�q�bW�a*"&��oڎ�sڕ�
�����{"���
�AL�}E4�dB4c4�`XNU˪t&�"El�0��7ҹ�����r���ⅸw���
��c�0Srֻ���/�v[�&:���>tP(ԑĐZT<b��N9<إ���R�c��7�׹r�%f�#�r|�K��B>�CBw:q���m�8Q�yvY�.��N�[J�4�vY+vѤ��-_���C_��t_�-�c�"�:X�D�@41|մ)>��O��^Ǽ��8�bU%G�,��jw����oۯ����^ 1ѽ������y`S������λ�
����QxM�sVz��� G�Fy4��4M����)K�)�H��,��Kf��@;�L��%�h�b4}�w�ŋ��L�,��">�[�I�����J�)���)��=�D��S���L��y�����G�mlqu{���m,�f���N�ɹ���.�}�O"/�-���r$��g��2ֈ��w>P���w�|�c>+.J��~Z����/p�2��%ΐD��X���d�]A�Pj�k�4�s1��hP=����]�[Yv�FGP�JU%��`.��Kkc��������o	_ j� X
�6��G�?U�êPV�P͊b:oO=O�պC��9�>y{��yz���!D��d2�L����j�r�r��"X���P��h��1�S�p��]|��|�JD=Ε�#E!�4�f����'���������{|���?�'����ō7�y�:u]�
f����O%ςǹD/
t�Ȣ�8·��������$�����R�|U��ǹ���:^���%�E����Z�5N���T}0\4��G�(E��$wp�uM�s�jʔbi�v�4���_����H��B���h2(��{T��)�#�bJI��[Y��**�f�)W�z���AEL%��=+]�	X�	�������5���g����=qV��ʤ����d�u����a�ڳ��jf�tB��Z��C<%��, )�.��HsT$'�4GJs�'�����U�Xl�������k|��B;�0�6�F����N�9*��`�(=Ɠ4\O��=O��]Tw!����=.j�q�b��|��'E_��T�=g�����]�d�T����Lܤ�⯕�~�CZk��%on�������{��?��Ye�nؾ��_���o[�/�/�#W��;'���ʪ�(�<�R/7gɥ����ޣ3d��q*�T0�f����r���ݻ���e5,j�J�����f_b��~l��p���*�{BLfǄ��5�;�־�˱�F�"1u��M�
�D�3��y�{���}�\Y�� "�F#����z�*��Cf����J�mp�u�l�Zvc�6ھq~�͜��ҷ����/�z�h:���z�o/r__��t\�M^,����p.�iJ�rb�U-�|!)kG1�4�Y%���龰�?p���h���߯Zw�?����R]��
@<f�qP�n�L�!K����c&���z��㜊�Unv�N��a�I�k��0<7�[��TW�1&�����$���x<��_�֭[E�d2�������5=Yr9�X$u��라9� �, �9>�����GL&ڕ��,����ƍ<������,J~1��H�����:���"��eH�E�E�_&Z�����/Z۷x_�h|�=X��oï��^�(��C�ab9%HNπz�	�D��Ĕ,&u]w��/Z5_�pD�/
k6�7����i|ݸ>
+��mU���B����[)���,��e��v��4������=Yg��91��/�y��L���HU�n��;�\�o ���5]�E��5��1���ƾV�eI�u������ܾ}���888���K���%���:	�D�����J�ZrTՀ��rxx�����'��+���:����F#�s�S��d��e�ȹek߂�<k���n�/�'���i��ߕ��|���1O�fa�\��"��R�w�K,����ɢE_�����M'|>p铨j�-K�$�Ɖ�WW>�����VnnŮ���V��;gj&�E�s�[�
�h�o;�,*�8�w✊����RS*����ߗw�yǿ��;�Qx�?</��
ZO�f�%M�S�^L��Y���U!����^	�0H��#+M�� �Rp�"�W���8�5�l��}dJ�njC���ʛ���K�)7ߒ	Ww����������x�QY�U�æ#T�(Ig�2�Ѯ�3\���-���:��G||?�ze���IG7����u�+N�#�UX��CB�����(��$�|͋6YT�(��&8�)6��QB��9ae4 !�.��Ɣ�*�2��]G�W�$�	)���dXה*��Z�%|YR�
N)�m�41�LH� BhI��f��Afm0��7D�1��x�D�xQ]�]�=B��GB	(�(f���U5�@�em�fm͑bK�[�V`]��(E�h��pP���`�����ONh�Hj]H!2�$���%�0�Zʲ����|�&|m����nѻ{W|o�}=M;��ܻ�y�ߚ����Q�v���� G�bN����<��L�E�'��FD"��E^T��� uG��w�ύh��&��P�[�-d+jjs�V�9��l��ǜ�R����I�eH��hF�Pf��b�!֟B��GBBp�ߵ�v}PB����Ғ!��G�C��1E�A]��<��N��
�\�H\��b�1:�m�B𑤑 "������.�,�GI��Hj$I�CA۶e	>��Dт.��%j�R��@U1͙�N��k�x�b��༼a���J©�Ԑ�0u6�4���F�릙+�L�a��o����{��J��6�\�t?|�*J�K����_����˓�ͦ��n��5�BKW���T�y2T���H1��D�{�-Ɖlau���9�'�6��>tz�ʊI�Z�|��W�ջԑ�������Gw���:��_^Hʖ�$�r�y���V�%��$�rF۹��Ia���R캆v�B`8T�j��W^e}m1��>��#&�-P4E����B�����4���ܿw��W�P;�Kc0������&m�f�'yB{��X��-/�c��J�B�������Q�pP�:�4����l�t2�x:cg�hF	\]Ǥ4M��guu���5��֩
�w��}�����g�]���.$�]������L�)"1�$e�Or�*/ζwV���b��9�$W����v���u}����eX�z��8:�Ӷ0���!����9�`�>�~�!~�v�?@D�q����ҮO ngD]EP[��G���;l���rf�,�>#������qQ�_tϟ���CDR�$���b��0�$ 2q��dFgж-��E�c� ER��cR���dK��"��9M�[pYV�1&F�F�Gj(j$�#.�G �tr�^�!��������m���yҢ���_�����'�X(Y�H��9�-�B�RD5"^Q�UE�HRC\n�$	R��8<"�� �)R���S
W���fGQ�"���=J)1�:,����:O��̗5���Ec��gfQ̢z�$1o�pH�vʣ*s�L�=t?����}a'���!��M�lX�8�9y�R��=[s�%<�<�,�$b����s"�D�j�hf)��߿.�o��{��?������GL��������eaQF���=v�>U�r)3�'�$�+�	0��d2���{�ܿ��X_�Yٹ�p���gv�p|<e2��"u]0K1[eW�z�	�D� "�63�����2�W���*+�5�_����[L�S���l9Gz���T,��\UYor��67�X�\�\gme��.k 1��89:���]>��3�|�9�Ʉ�:,��Jԕ���1�p��k���k�z�ò�,�{ۗ�h��+�)���@�6��������������w�����w��	�,���O�(��V�^L��Kp����-����[ߺ�͗6Y]U,uЖ�d:�<��Ǭ���o����xX�K'�����9���h�"ބz�M����H�^�Ef�D���8=	����蟉�2AL=�9�0�����:�D�[E���\Љ��D/ƗɞWn	���l���?��	ƫ�|��
������&���J�D��t��p�Zb�������r*�̄����5������e�C�D4!�e�-9�f�)[��`���Y-%0��zo�|!����f*�rZ&�����4�u��Ήa* ��G��>�g/�W���p���DOz�]�L1��s��O���m�SB8ˉ��@"�U]`�ֻe߳����8�""�Du&��P��+dg>E�೎/���ƻ��������_�8�MD$���3U��~���X�N�I$��&̒8����Ԉ9�yդ�h2�����:�o�?z��O�n��Ē�9AΖ�_�b՜�(5�I�G���ߣ�;��"tDli��(|�O&G|��8_҄�nMp~���5��<b��>'�S&��m�fWMO��'}Q<N��f)[v��޿�gkk\���K;#�;W_��˯p��}��'��UD����b�]��k�����׾�[o���[��X��RQy�I�*
�ʓB�l�p���hQrr<a:��R���Q��Q�%W��������;�e{c�A�
ɒm���J�D��хDg�:������m�{�3>�U��;w�����s�e��E�w�U*��>U��A��p�[7_�;����z�����)6İJU�����.
?�iM���g<Nܺ�&��X[����s>��
'�m�	�*N ��}A�	�ق�-89�֩����I�)���]�w6񞒼Ǻ̗�\�*zRG�\m�@�X�/�u�ؿgbɤNL!H��M:{�Eu�t}�29���"!�P'x)p^Q�ݜ�v����]����M|?��߱�6_�إ����1g�i�3�xvOK�{9�5d]G" >���؞�W�!����Tɦ�6Sn�9��Ϸ�'��9���{�$/`�?�GWdKe"��ĮG#�@��|%�-��BL	'�� a��.y�5�O�ED��&��,!Qi���Hw�n��YbE��1�����:�Ǣ�vU�C�}pN������2@_����Bԩ�:ˉ���W�G���.�|�0�K�EM��>g3�#Q����$�ߥŔ�����8=���σ!�pb4�)w�|B�ɢ(����aUS�6ؾ�
/�v�|�§qxrHA�a[�i4��EOnP�	��|:a����L�W�յ-��t���)�=d�Ͳ�/٩��qH)���S��<U�,K���x�����w�ŭ��3('���$u���']���������](IB�y��5������׹v�5���Qj�e�DBgFH�������kEQ��oP���ؠ��/����R�k�Ǔ-��5����^ӂ�H�=�p��K��\���t�	�k�h�������6��P-UA:
/x�Yۺ�`4�HI���=�yC"���;�uH!���N?�O�-2�ҩ<�{.+٪y���Gc���v��[-��M�������!�d�����uvCg��ٓ,��P�:��@�ԏ1[�]�O�ʧ&QA{k�j&��소)[������W�=�_\vz�2Ձw�ښR"Z������T��-�Kz�Z"�EW��j-���RB,��e)e�j2�E�1eˍ�C]�J&X�Zx::��� �9!u${H2�Σa�A+h�Ę�EYP��y�h�/�+=E�yAd)�6�4�K�b��H�w2>��-0���߈�L͂!��ⱘ��W�Y-���o���i��&bD$?7jΝe]83�\���4]�Vg�R����{s��z/�S�n�0uw�|c\��x1e�4&�E fk��<��w�pI��+l!8�~�]ly���3I��C������b2f�������JO��-v6j�шՍk�|�!v��m�MNH*$K��\����(��YJ��b��落�����2�`<������5��'Nf�E�.,��E�Lr{g��pu�j��jM#Ncv�i��󖮝�4{w9>>f��h�&뵊Q��($E9b0�`P���D-�fmG;��t%X�F�o�h��y��0ZYa0,����2�]��|���!���]�/9\|��Mx0���b�e�/kB�bN�ݵ����>L�S��GH���56�����Wj�VG���
�+�ll�ě������O~�t:�=>A,�4�-N-����
��ɹ���'�D>�@��h�x�כ�Xv���]Om5���GJ�.�g��D9d8K�9uX�P�M�Z.����s�E�Qu�k˚y����8�p�'���2��|�!e͞�~��k?S�:����ړ��I2���B,I�X���%�1�]��%��^��\~&GÚ��eRo �Q�\ͧ���-s��U=��=U�y���L�9��	M�е-��u�)����*����>k�����*!VV�X[[��+��$��	M;gz��.[lEN�/�Ӭ}Y�����a�H�%K!�4 �˔$�nv�8�pxX��;u�b�*`�K�_�a�["~}�?5�EQJYV� a�N�N4�>��?|x�)N�K���H��۷=쓒&g��Ÿ���a<�l�[rS�Z��K�I�)�)i3��D�J��a�if�ܻ�	X Ԟ�^��+׮1v��q	��f�C����H@�1��h��I!`��"�9��c������\�2��W�X��a�����C��%�S�ڴ7H��d�G�ޣ��̚�q]��1`\WĶ�d:c���}~�{w�ppp������ߧm��Ρ�A���pEEQV��6U�5S��vyp�{�G4�zw�pr�G�Z�j0b��^�z���V�ͭ���C�2�n&�y�|��FL�l_��hD{7�"�	`JB� ���p��>�����    IDAT�����|�*eI=2����ڕm�]������!��*W���`��������1��N^Յ�,��Y6'8�42TD���)U�yr������%F��E�ʙ'HUz헜Z�R���αUQa���"��k�򂤯� �KS��Q�1s��(}EU8W�
Ż�d�')v�d���ު���j�Eژ�UU�����0��c ����5�vJhbꭔ�E�`KOZ�wc��Ĥ9��N��/D���^�[��VB����sTUE]E��8<4��	)�)�(r_Ԓ.u�%k�o�2���w����l����|�	��1 �0R�'�]��<�������+�5��ܽ��'�E�h8fc�7n������늢�E&�C����}��qpp�H"���/�%W�!j�,�!�R�
# �Q�>~&^�Ǉ� IUI4�L>�"`@]�Rץ��Z#!&	M(�s�{��B1��i[�Yx.�W׵��t�%"9�o������:��{g��lh_�J�'61��B�@�k"Ė���Ķ�XK,
��`m��z����:x���]<���fKR#Y�cy�.��L:,�ل��#hژ����5�zؓ�D�F��vq��u�#n^��:NNN���A�uL�'ܸ����q�����������_���l�rT�s�e���W�!�+�,�e�#�4͌�Ç|����/~�ǟ��d��FO2!t]H���V7���-fM�q�Ǭ�\y���s��O��ϘL���~���ˡ'B�~�(&S�	E&$�&����?�o�����ܶs���yO{��+�U�W�\�Wn����o����:�(hlll0��S5���XZL��w��&�����}x�4��ʗ��_�,t�
KZP�>PDZI�������G�ѣi�k�"!5���Ɩ�����ら�~�>��f���ˬ�����J=P�5E]�R�ifL&�̧��9�����v6��|]�Țؔ���pȵk7x������u�
];ez|���}��a��=��t˜�}!	E֪�Հ��-����rt����=fwwYT�[�Bz�bo&	⠨+VWW������:+�1�~����9��4�H����Sams���|���x��ׯ1��������)���D��'|��'�u�g�9xpb�R���Ң�%h�˯���o��������&�̻@UUl�o�g�����op���S���ݽǝ�?�����l����%s9���pj� Щ���If��c��I���������P\��E�W"-{���A~9�i`�eY�`P�JS�� A�%)���mu���7���e��o������ruSuE,�I2Ra�Y�{1�	�����V��}.D� �]?�)�T��Cb_%aq�G��	]B�H$�w$1b�'���=>��R�z�7^c}|���d��u^y�u������4�)�ù�^����;ʅ�.JW`��	��s%��p��ع������.,�G���<t���eA��u]����;�;����w�bu�fex��h:���G1�Lr����X�R4[L4".��������T>���~�7��_��g��bT4���E�1A�2k#�.��p���m��/��@�������6e�畓�%C�z��/�<a���E BE�T���b8K�4�l�U�"t�޷��<� �I@H���!U5�ƭ[4m��kTU}Z?x:� �SV�m�z�TՀ��b42��ٺ��;9��,�I1�5-��CN���6R����1u=d8Z���fY]]�I�C�����u���(KO]ק�O�L�\��V�ϧt�c�������9:�2�wT��s�S/��W7����3^Y����6k�EAQUT��tQb����{����������î��ҧ{	8�qEE�����o�������IUK��h���}����w�����#U`���D|r���Y�R�cF+�������}���u>��~�ӿ㓓�e���^K�������tμm�Z�d��	�x������笭���l�K&�����pER-!� _���ş���?���q��k+���ks��<m2�YIkc��dkm�O~3��_���kW��!�9�lmo�}�*߽�=��G��@�[7o��+o�֛�amm����ϧ$K�c���Nloƽ{�N����B��������kO4V��;��73�RR����peݚ;��O�#N��$���"2J$ĬO1d��sc�Rt�-��>P�(�Sw$VV%1F��EYX5���j!]�X��R�?wItu�&���[�_'���omŭ�s1r,$�&/�b�­)�q�.+�-m�xߧ49WbLU)ʬ�S���LC�!D�)�n���]�ݽ�����J�)c�\��ε�q���w������k��EB��}^��m98�P��A�+��U9���������a��:����	����f�>�ri� X�t��]/\��f'�A��d�1ϑ�d+'��&�Z2��f8'�pr2���8Ga�� ��8�ݯf����b�{�hh(���Y��3(+�Fe�ꜘ:��J������c2mh�H4��թ�T]q�7��M@�*����֭[\�v���uU}J@;�m|�O��g�?|�g���?c�y��!Z��$aD�V��4������6���:o��W�]cu<ƕIF��S�8��8�EQK̛Yւ����|���_�ɤ��<�/36Gk���k���M�������M����w�:e��x}���Y������ۇ�g�~�����LF�x���Y]]gck���+�olc�cPy��ʠbmu���;|���3�?�Pl�p�hA=�}�*W�^ge}L�"&�ٝ;4M�l�҂�(]�D��`D#�a.��������7YPU>����8�/*:�62�޹���w����׮]a4�4G)�FN=Ml��A<�H�x_CK��-��1{{{Lf-]�9Q��(����D5!�`gg��������_ccm��x��`p��s��Bb6k������=<x�l6���RP��=B���9<�=�>I�)Q3Įn�)�������D����%�8,X���{���B�^��x�$X����������Xx.����8��z3�s�d�l�=z�B�Xʶ�b�E�OK��s[�؄>|��L�'���w5����m6��E�0���]�T5�w�re{�c��Wo��ko�M��p���r`h�R�H�esz��R�tm�d2co����u����YY�dee��f�<�i�����?K�v�09f�	]�S�(r�F\��,��J��>��"@f�,fk\�!��9E��IR������0U���9�MV���˝	����>)j�OA���m$�
�E'BUЀ����� ���,P�!A9j���n��bEYgW�z\�H��h��ԣ1/]���[����os����1������)*_P�R��5�?����
��_����M�����,K�	]H�6ulllp�O�!���?���k�WWr MO2���hq'�z�Eb&{Zd�_j�>8��;�?�Q�
Qq����������z��ׯ�V��AY�Y��5�����@�P�UΏ�uY�N�'��1kZR��S�E���\I��J|5ė�a-lloQ���J�H��u�����mmg��pŀ���y��^��͟���>����R"'=�jf�[;W��wn��[o������~N�3�mnRWbA�r�:߾������W+����4��n��`�(|��y0�:���à�p���������w$s�j�p��xe_V����ޛ,Ir�{~�����1�\��YP @�H^ކ�Lm��`2�B�2Ӫ��3�7��� Z���nKj�� 1՜U��c����8�Y ,Ҭ/�VȪ�ʨH�����N@������p5�V�f:�q9>g>�3[L������S���9:<d>��&	�+N(�p�����^|���/�&(��@Q�����F�sA��������fK�UD��?�m�d�t%:{���xM�<M��tF��s���?O"�v>x�%D|�����*>L��cR�VN��hV1cK�)�=�,��V+�F%,���"6��!K���S�>{-M�;l�;����orvz���*;�#|3~v,��%(DB������t�x��zA�������3jy�?^m��Bo�$��Z΢%�j��뢁��W�|�3K��	��4��� TD���_�Q:�(
�}E���01�!"E�1�g9��+���sͺ��cV����ݨ�B��`��G�C�h�Ӡ�@3&N�,�hM%e]T�QXg��C������;��g��{����W�$x�AI�.��J�f]R�t�nT��NN��0��	(6Z�8�ع�������Oʭ[�h��qL��ZTW�e�"��*�����y�m���ҜCh�r666����w�{�t;�L'E9ie�d�@����0��&K���cgw������\�ˁjQp|z���S���n>���bI��	���k�7TQb�H]+F�9/�/xyrI�u�i������f|9����$1	N��l�D�w��sc��wﰾ��N.��x��K�|���d�B������~�.?�����Z#�R��1GϞr���ň�d�
�BJ�N��dlo�����v6�v��Zo"����fT�RV�����m����~v��z�Y��G����.·L���sF��XE��u��h⬢��O��6]>x-!hq.!H&>t�"7e9��*F?��]�e��e�Y+"b�^y��Kſ���8�Hh솔x	`*�&I^�ܿ��q|�굚�>@AD�	Nh8z�b�����"?��	��&x�m2��5n�챾��.�39=?c>�7#�f�1�V�4����G]MPi�+�<���`���M��6F��m�`��.k�,�b��"7M$��Jc���j泂�tJU
�Q^����������������;�5b�	H�����"c_Or�з�(^V�[E����AB�QT��]���a��G<7(�����a�U;*�s \5�A��A_wQ[5{+�«|��	�ST�F���o+TH1>ڸ�(�A!J�Zy�]���/�.D/�X_�tk�y�������O�m��tp�1��#+���<��ՖD<y�IT���]2��B�E���Ԉ(�����M�~�m~��coo�$m�<,���((˘kt�2:v.`m�s��� �=E9���)O�1�W�J�N����m~����p���<�[Ǽ�y����/�/Jfe�d:��6������:[k=�ַ��V֎���E��
���C|������s��m޸u��A�4Mpa�kT�:��ʯ���WY�$�*���������F> Q���7�����gO(�K��x�#-��������oqcg�V�x...��g_���Cfe�$)e��������wٺ�K�Ip����#>��#?���b�eP��E�v�s{A7ﰵ> ��d-���-�V�Ӌ�_L�$E'm���JR�����ذ-�~������x����,��]��ua��F�%\����~���+|P��H�}Ȕ�\�M�����^zý����s�1~s�ר�\PF<�;'�YQ>i��פ<
(�F7�R���9�	���^_��TP�뵚�?$��/!(V)�MW�'�RE��d���$��u����޽�9ؿ�5�lcΚ,ϥ���J�"�6�F�z�I4�\^����s�n��9�y��.�7vٽ��d6���"*� �K��=7��F�9�x�f��|��)K��G�}fV��W�=V��`S|��-1.N9נs��)�N^N��h��􂁠�C�i�+4����o!�����S�h�5`b�%����EX]^"�P��B�Oy�Z2
\G����H�!&�xoѾ��̅U��M�A��R�G�ΗjL"�VT����=���n߹�;����?a{g�f�(8?�����dBQU�pɀDJ-%��Zl���S:���5(ɘL+T��%�"ow�qc���Gܻw�[wn�j�(���s�<y³g�h�q�S���c�FJ���0"ת�*g\^�svvJQ�h��TB��r��]�}�]���0F���>~ʃGOx��)�Y��(~Q�!�s>�����ҷ�e}='5�4'��D��z���r6gV��rR��]ƣ)�6t;��[x7����ٯp������QB*��$����鈧O�s��.���5�7n�`gs��ጲ��������g��-�N��Y�1Ϗ^���3Ƴ)"-L�Q����6���(C�e�ł�|�pt�x<��/�֓jSq��͠$E�%	"qj��t�����$AJ�$ }v\U�责���9Ϟ<�7��/��8?��\�DE�e���_	/�(�ҳO�`��Q�r�$@)&���BK���y�4|���������g�uxSB���T���[׫�;����%oP%���]Mx��y��������՟��o�X�U&��"�mފ���ky�};�@�]
I${�6��=�֝7IjO+����9NN���8�]fs�k\�
� �����.�y������t�~+es{���999�r4k"IT�͸48$�h�؆=���WYYL&��666�ی�l5Z��(B@y�8�wq̫��#K%t�E$o9b��d(�QhІ�5�ML%E�+t�1LC�F�(�p��Z�H���c��X>D���x���T���W��Wk�<{oc�l��iE�j44���Mu#U1��	E����}��N��`ݜ�Ι/�+��N��������7�bgg�0Ox��9�>���!�јEY`��J6i���@;��{ܻ{���8������9��r�r�hz���͍=~�����~���&y�CUU���~�'���/�#?N����^�ٲn-A�E�ź"�D(Eb4i�����ݻw�qc�ԤX[2�y��1���o9?��|8�v�J[�$A����rD��T6���(���;��+vw�9::��!�@e�x�,j�(n�9�n���D|��Y�_���vH��S��-J�>;"o���;wnq�(v�6������sܼ���0�����}�.7n�@)�t:����|��!�ć�R�� �£Y�Y�{T�o����u�EE(�.M��J���.��798�.����k��D�Ơ���^���΋�>��3~�O����e�yZk�jb݂��]D�}�R�%�k���Z�|[�_w�^{���/���������^6�E�w]e�%H��36ت���X�&K�5��^�h��"���weY�,�V糿�_a�V���tU�:���!z25{�׭���"r��-���`+��Ds~~Ni����Ռ3�`�k�3��(899���)7�{��B��g}s�v;�����j���EH�kޛ֚n�e0�n�ɲ
V�󧨝�|�����B�DH3���z帮>Ռ�B]⛍xxu-��T�Z�(�5X,�ɳ�,K�=�wx�_�����4�n���:_�[>���+�}�k4�$IP!E� ���eFŪ��"tZѤygg���I�YLLg��`��veZnܸ��FDe�G#NNN��ˇ|�駼<:�(
M㥄D�[T��7�����I�#������ޣ�������u�oq�����s���!_|����o9>>FI�l6��Dl���k�)� ����(M��F���^o����v�I���(T���;��Jst�"���9\dI��������&Y#ִJH�k�.F�h���T��J�e�0�/��x��$�#׎�/� �C�L����#=z�����ۨ��	,��^�h��H I2n޼������Q�G�<?<�ɓ'�F#�fZ�(W!:'5i<�"d�6���vsnݺ�Z��%T;��THL�H����kl�]P��H��,Kʲ�A�a�>�G������?棏>�W��Z�h�$*6˸FTuu�,�����]nb���J]�}��u��\KgfM�j������?���~���l�,���[�[7��eL�s�y��^[k��R1Z��t����c�EI\�B��q��R������_|o����z���������tT��G��d    IDAT@�I|���U}�y<�D(M��d�+$�A�����{�TSy�A���Kϋa�f�v�O��ؿ݂`p��#&�)B Q.�?��P�p��ʕx*��0ڒ�0yn8��2�z�<퓦��1;���'�Fl��Ȥ�� m@��.���8&P1] Ҧ.=n1`~vJ���*����7�7�}��W�4�8yV�! ��X�9�c��5�h敥P�"i3��VL�/E�	5$���zM A����$x3��'̫�m��.yk�v��1��$9b��9���.�g]t�&iwy��>?xs�SB&T��8�dt�sbk��Z}���]�-y�|�� ���)Y_vY�gԕèA2D���y}�!z��,���1��8���}�;�w�ug@^ըI�0�����?>���(�i�&�A޿C�o3�Πq�����f ��{9�BSzK��RL`kA��|���޾s��~�j���x�%-��Zz���_�	�������cfG��я��Q��U�����W�@�v !���s�Jpd��&twY�%-�T����������wz�䴶Zm�4�5&�X[[�;H�zG�JQ�9N��.u�#oH�-.��O���EB�:�qA�w0e����N�Q!�,>�H�ٿR;��P8�(��C�R-9E�K�82���n�c��/����_�O��O�͵�}�m�j��=Ϟ>�w�����o�霾�(U�I�p
�n�kn�z�����,ׄv�{Xզv��VD�Eb���yYF��Ω�0�O)JC�Y=��s��>�!e��nVq���|��#g���}����3pe�$!*�E"��-��K���ٔ)UƽbPT.�i�`�ޢʂ��V�٤���R���myO��>�M6�zk4�%�0J����x����$�������� !�R_-P�N���D7ݸ`�f2�V��I�N�T��i����4�*����� U��{��T�uJ�%(�q�k߿��������^W���$+h����9��e��O���t�pt�h|�V�&1	��W3���G�e�t6n��$�¶���D��2�]`�������s���m�ӡ���v�S��q�k
~����*&�	��^n�TV����Q��^�}W���6O!�t��F�h��"o�ź&p]��,gms��7�*��P������Y	*�;�`��>o������Z	�.�8;�уǜ��,\�����ӝ���r��E���������{�E�t2a:�b��V����N��Fb2��n�fkg���-�<��/>��,�9���DY��Zk>��i���W�]�VƬ��,� hu2���mm���esm�^/��G��GF�	T�bQ-�\����ǰ����������y����B'h�%x��ټij��ڤ�A$���N�,	�vމ\HJL3FLp��IIL���Q%"c��Xg��1q&X��K�窕�,ƀ�
������چR�w��MC|��m�}�Ngc���8�ء�f�6�޽���g'����޽��۷����9���<�����,3D��K���@�V*���	�3�qd49�$��qA���yJ��Z�V�6B��|��%'''��q)�h�]���0�8::����1���V*+����{��4Z�$�։�i���A1��c��p�>��? >\������'y]�����n���@��R]�	ޛW����4��5;�oqz�#z�d��6P"�9+���?��?������������z�����3���6!��	���Ңoy �dCp� �<�W�'�����숃�,���2�Q�)����%��S-ב��E�ƍW)�
,�.	v�h4�����l�n7#�r��y��HL����(_�����������׻��j"ˢ9��5}���w��B|��k�RB�bk"�|=.*,sa�HX5�}�E��e(T��������`0��>�$�h�|^0��=�[�tY�3N�^������׿��0�s-�$y��t��W�p����4N��K�B`<q||L9_0�ssw��`��"{�>y���pȳg_������?���xF�b�%(�,���'�s�v�fk�O���LB��1��'hI1�Kj$�Ҿd^�Iۊ�{�p$1^,$i	�|���QQv�iuԊ?i��:��<ĦPC��$���h�)Y��q�uAK�vY`�����Zu�u��^�H�;��c��Z.�%''_<cVN����j�Ij���I�ZX7���ԾB%�nhiH&1�f�p.�DΝw5"	���
.��8|򄃭���5�z=v�n���?"Ks�o޻���-��.�ل�O����CF�<Y�!1�9*a%f��`�!���5\ښ��S,&T�ʥX��ϑ���xo�
噌/9:~��'O8|�yQ�t�h)-��4���j�q�"�R�R�D�\������%�����u�*��	^��D�J�ȮJÖ��y�ˤ����{z���/~��W����?���h<>Ͳl]'��^!��#ڈ��Z�e�Ue)W}KaLs���t���M�r��~��1A+%Ai��!�F��y"a������TR��u͙������IxM�
�L��S���b@y�R��huKUL�O9?;b:�E�B+�HҢ��dk{���\�_4Q4�@�W�I�o0~�1pVJ!A��QU%�٘�x��fT>.5��.�:�+b��9�@Y����7�����Ѷ�Ղ��A}Q�xƇ_��ӫfԣ�Ҝ:D�x��(E����(e�Q:�3X�~���]�I	�Py!1-*;DDa�6MB�縺b:�ɯ������3f��		����_v��I�1QMmd*D�V�E��A)E�=�E���;;[�Y4^���(�Ŕ'�>��ɣ�py�t/��/:`�x(}�����,�2	)�)tPh��i�D�_'�x^N��iQ2��)�%$����c�b�Qe�!(�.T��:�o�77����`Xb@�53�f�Dى�%&r�$P�|(�PTT�)ò��:z����U�s��ZB������ٳ'�������!H�&�A)A)�ҁ@���2~t�6��B䲪&�'���ޡ�4"�D�S#xWq9<�<}��v�[Z�6��?��w��更RE����b��/x��g�'8_�[,:�x/,=���F録X0:�����O�YR��-XrjU������+�j����t���H�I�ީ�z��cV�E]a�IB]�WԐk�kR�^����υ Uei�rc�$A$/-A��}���L�<TU!�^O��n����A���T��dY'�z��ӿ�ȏ�u��%�:S�eVV���9|Ղ���WH�7Mv�
lcB�""��
<����+k��V\��9��#>D�Y\c�-#iUK�7�݈`�EU$�;�lz���s��ȩm�h�!o����e}�����$����z����2���_�o=x�r�p8d:��� cZY�~-�"B�jJ^ݑ}��s�f��`���L��n��x3/�?p̖���j�7:�t���л�T� �HZ5i\�y�j��q$�$	:i��Qdy�v�M���jaV�(�Ap$IF���:PU5*8�/Ny��3~������)�t�Q	�����I�&��x���hcل(Qe"�Iw)��bX�ɑ��W�`H�൥���Gǃ�e<<"O*
���:��FH�xm�����<Ƥey�Ea)m�V��m��*�(�0Z#�B�cr9���/N^2�Ϩ�8*&Մ��2:4�Fŉ!����
���� <4~E�6�RsM�(��@��D�T@+��btq���Ng#��Z���sM+���|�t:���X׎����.�gq�e""�Q�DB�Fi�I&�
:U�<���m�����I@�L�J�&<�q�W�gCN���O;dY4��Z9k[�l-��������/���Ǐ2��"(�ƈ�#^����
���E��<!K�Mk����G����C&�&ic���lؠe	Ҩ��5����(�bm I�>>Ьe��kJ^��*'4������Z��U�A�އ�u��e�
��
��V�8��7?�:yxy�8__�닋Too�rx����;Q�����!�j�8rJ����[�B?�1ʹ�Tu�TUi����s��2h��
��jσ��}���B*Jk��VB�j�oz����^��Õ[� ދ���-[�W�9ML�pED�DS,.99~�'�0��x7�t����8�h��u��J��l���q�4&����i���l��Y�,[tL M���}�,g6/vD�b�ثuݪ�V�D��׵t�ո:6�ZA�#��}�`�J�-V#��AGT��f�7F�e9�Ic"��h>�tT�zE�^%�i�Uѧn��c�(�1:?�����GϢ��GR!z6�i�1�n���5Ƭ·J���ʢ����GO����$o�u7��v�R�Ep5�ٔ��3F���bM�C�9�I��k�$(�N���삗����<!�:EEQV�N(B75>AH��_I��H�x����_~���h�i8<�S|0(�V�N�G��f:)�6�/�ll��1㎈���(Y��b���hţ���|��ƀ��aK��hƳ�S>z�%�ш�l�B˽�C�A\U�r�{�L&��c:u�%��(<u��h�:�IS�iP~H[1%o{��x[�G�(ݼ���K�; ʡ�`�soy���wYT���$�:�
X�N��t���S��O�m��$��x����@�%�ɬ�U[�<#1m���*t+mI�
	<8���_c&�u�B�����l�٘]�VYnڜ�]կ.�W��oF����~��)x��DEDi�m0�����|��ϊb2�v����)��]z
���� ����4�x<֭��ot�_b+%::ŖE��L��^�#�-���"�z�[���h���XV�l�F�Ң�(Z���������^��+ct��]�Ba��-�4I�}�%M<��-0J�U��&��{F8Y��JS��M�6�������./��!�$��ɑƻ,6A��Ҟ�.���C��Nא�ڬ�Ek��0�̿
��~�k�f_�����ﵓ�G�xdV{s���+�/���j�_q��o�b�4#����)�ݖjN�5&��Яb-�ق�dĢ���5��k������������UE1��'��Z��ʤ�������fιՃX)MՂ�d���3�=����q9��]ۤ�
k���HM 5B�
�!k����`�ńZ"oL�mZ������
cbsrt���G̋���'B��D�^C#
%��L8*.�#�ʣ��Y���xhe	��wnߣ\�9>z���|5&�bJP0���L���a\�XB��傋�S��Oh�����o�L�V{�2�sqq��:��@ek���.P���
-�o�˫H���1'8�b�b�=`k{���]���i��Q����7�X,JNG�J�5�]�������z�x�s�P3��<;z���ǤiJ���h�jŕ����%�|F���q{�F8��F�6F�b��b����t�$�ps���t}.//լ&���;�6�t<f2�dQ�i���-���=K�]fl+uM��$�HC�_�ZYZ.5�_���⻖������	��|���S�|��I��Å�^�?6J��'������f#�pz�~���?��������1���E9wO�q�*+ŢJ�"��f�?���V����^9Y_�u7�Ʒ�9PJ��*4���('���̿���^/��T$	�DB��κ?jIY����Z�W$H��ؼ)#TuE1��=�����z��\#��m�����B�eE$�/я@l�L"�V#���Y�I�����A��g|6�[�v_�.���\��;-2�F�\�7�^V�+���b���D�E�Z,V��Չ�ʸ+�4&�:o�����(�'g'<{���'���1I���6n����{�9I kKL�$&gmm���5���UAY.�E� 6�������r�~}��\�x4���!���>���#�<IQy��;�c�bVVܹu�!K2Zy���Lo����EM�
�3L�ct�w��t�W�,�X__����z���K\ KeI��rV���x����.��%Y�C�d*!x(��ɘb:a1_���Nw���w)���Ֆ�\D�OPH0� ѓ0�wK�P�ӨA�;|1'(�r���/��i�LF������~�ڠ�˗9���6 UUD��tJY,"�aqδ���B+R�!h�7qC����&a���`�?���w�����bm}��o���t(?{@�X0����b��2"�w�v兠^�<�����no���Gy��f��<}�gϞqzz�W+iL��xo���q5*Tԕ0�sv|D'KI�gm�����n��[��ՆO�Q	Jiʲ���'O�����OYT��}�Fk� ��gt�ED_�&����B��Y2z_��yK�Jϑ�D�jU�E)��4�`���Y��cv,�0׋4mϒ3��(Z�V�_tC��{�%�On'm��u���d���Jkkq��lj�Z�(^�̷��~�K�~NW�h_�zq)Q!���Q*�J�|��߿/�����>��C�I](iϕR����ת�-�j!J"�D�х�
ثrt������j���>�B������^��;o��BQY��6��������S�D���$11!�l�Ѝ���c]�u���
7&��h�������6�OO(��t5޽�9Tl,E�>ٲ���ż&�ID�p�nB]�e�FQ7�Ө��RW.B�ί�4�4���\g�'-kG߾łn�����[c2�EkMh�8�[!r�.U`y;糇���������i4���<~��gsn�Ϩ����M�Y���N��O~�3����#·�r��Rʪ��KT�"�߾��![�&f��g�����j���)UU�����������W�LQ:�פY�|1���2^�xy�_Wܺy�V�!o��w~��`���]l��	E�qV��Z^�8���%7����	���m����4>��cF���b<�ɵCD�%Q!�g>�1�Ϩ���ʨm���ʒIF��|��G�����"�Ak���]�Ii�Z�L��s�kOYG��[$IF�g-�
WVL�#./ǔ��	�����c:t;�l��i%}���u�w眃��eI1�9�g5u]3���8���ϟqyYPۈ�4A����
��߿�_������{j��1�� ��ǻ��=�{���7�կ~�d2i���,��6E���,퉪x�7�[G�Փ'O��w�~7��2�jA����?��������@�c��JҨ�vok���G_|�txNU��[?�����N�v7G�h���Z%X�wn����V���c �G���ʹ�Y[�S�\m)˒�dL&��ycU��i9Y5����7ڱ\kJD�r�p8H҄�*�i��I˪hk�Z���5�����>�&�����Lc��A-���i��m�~�ӟw������mv���o���m�H-BR,����$�$"�����<ֹ�O�r��r�B4�.�Y�IL��:��H�D��!��K�����A��������㏿w�(��z��������T.B�^��JI���?�u��fÑ�*�X��=k|�[TH��cU���/�NRҴ�Z��HCr��6�*ߠ�}�_I�Ccyʲ1�C�q_�7�k-��R�S�Yކ�xl�ڴ�4o�e-"v��[]Z�i�am�1M$MS�xW��BՃ�B�f��|�d:b23�M(�cQ�S&�F�3��9�op��>�kk�SC��S�9�]0�g\��P�|�Jd��e�z�*5�?G�j<:���R[����{��6F<�d�~+gmm�v�cm@K�����zLU9jU1�8=>�r�&��6F)��6*l��[���	'g'���,���"�2�&�b2����K����F�}7v;J���3��x���G_0�[���u�t6i�Z�:]n޼I]͗S���#ht-w*q�y(�)Ǉ��򋇼8���<�W�e���×t�5�Ulml��{��ݽRH���*`m��5E1g6��P��Fc�HL	���J`�����wx덷�ٹ� I ��*xt����l@Q�x�����1�$|��M�5/����?3C�    IDAT|Nϼ,�ᐧO���ssg�b>���Grޠ|W��cL��Fm⫨.����kz����~/GT�(A��zO�bڈ�)�^�;N���H���+[��<*(���Ղ�t�h8$	�Ʉ�(V����=4��_�{�[}�9ޞ�m�(z�H�E�:WՠL��R�?-�������ԡ���N�]�>F���_\Cr���W�ͺ��I�2���j�V�.�^��)�t>����|Y�}=��g�sN���!��c��ޙN�-����Q�V�7�L$s�
�t$!.N7��*s�ܽ:�kIĂ�Z��o�# ����j]W3��V��@i�E�м�u�Ĳ�[�dF���I�������[��{Z5�ߡ\"��g.���G����vz��t:=�2XOK�u�.��-0]p92�Wxp!�s���F���h�2��m��(3\]���Qc뀳0�O(&c��PԴ����f���O���NY�������PB���},����$^�Sj��[��hmQ8_���Y�!��;�yA�:X�F�w�X����[@r��X�̊9��/.y��1k�d�a{��w3L����6;��<9|F���5���V��D4x6���S~�ϖ��W�	*$�ה��U��&��D��cs�M;���ln�@�a�\|�/G�"8-�U��P-x<�3�L8�Q5�ʨl��r�cP�������Q{{�dgR7�  8D*���m��6�8����J�A��"��i]�L��)�����;�i����zl7mJI�C�Ao�v��{�#%(cb���jWOh�J������|N��{����?��'0	�c����L"��9�&x��������g|�EME�7����u�t�,n]���b��H���999c8���
.
��5���������+馚Ǐs9R�q�-J}M+4^�&�Z!P�:ˀs%!h���u%J%�uκP�Y�1E�MI����i˟�I=i-.��M��+���?��%�������� -R�VR�O*�[��&I0FW�z]����t��u܈E:�%Ѳ)�_˧��oЬx���9P[+�7����%"�ޫ���߿>��ÿ���[��W���E!�Vˇ��b��I{���X��~�<���k-�%��ɞA��h�8tX����$�J0є��W��#������o���1�
)�}u�DZ7���t^7On�Zln�q��>w�q�{��khӂԢ�܂��\pt��O�����c���]��ǋF���$�	��5�h���e�b4$ʠ�`E�XB5c|�ç�v�`n�ڦ�O�m�r�U��x����!����.OrdYz���{�="2	$�B�����j>�j(3Y%�43iQZHF3��h-�?@f�ϖ�^i%�dM�E�#gĚ~Uw=�F&����p����u�G"�LTݨ�<f�gDFzxx�����|�;8'�Z��y��:�+:���@Dh����.��k"�8�()5�Fxx�KJQ�F��-n�{��[(F��o]��u< �Y��Φܻw���h@�{k.R9a0\gta��I��̳u�*o]����y�i.)K���+b�kc:K�-�R
���p�.E��2k��oq���
�A�\p$.WxӷcK��V\�T%��P�%B64vE�,m��'O1�[��1��1���[����1���ѣ) 8�S�x��)�qC�b��� ii���*�f;����vΚ��T�6�͘��5����_��3��w>�l(�X4�o�\K�r�d�	 N"F[�i���	�4���G����翡��	��5�!�c���QV{�RX	4��wwB�3&�k�qy��!%�@�az8�����i޿˝�>��'�ۨ�
Vrߑf�!���/�~|��Qvw�u~�)W�΋7�n��@]f���y�����2x/�HmLM(lBJo��?j��vY5>5F+�ݵ����O�d�>�� >�����O���G:�����b���+�;�Ժ�lTIM3[�����d��nE��ub!ʏ�Ʌ��҅1�X�R��K�����U����fę@߭���(�h�h��4�XPe���x_�j�[��v	����:hD�JT$!��p.d]�vI�>��ٿ*3�9��e��-�MSVD�$��������2�_ЍkG�
���tU�!d�6�r�*7?��?���~��K��k����^�����m��u��K�؟Ly�7f'9M���p���:��m�>��|;����fF�5��A�jIi��<݆_H��#޻u��Kk�oq��m.]��<��g���K��|��[�M�Svww���c<x���>I��o�BR�U�%�{;�'f��{4�6��������}b�`�$ib|���/͔0�0���֥.\X�	��X���amT��ŷ-�ㆺ�D1�u8[`m�e���0Fi��w�&�;�Ƿ��w�z�2��̩z'�2�qX!j������u���N�o����SNժ�t̠OS<!Lr���{̏��b�!�������*�������|��`>*>v��C��Aei�	�}�k'�lm] Ě�3��g�lS0*���'��<�������,")֮��F�O�9/A�$�~q����}�t����Z�!�-P�`M�B,��<%E4`D�.���1�����1���s�chĄzU��[bPJ��g:�#�Y��I$��ɴ��G�-�l���s������b�S8���Ң�������=Lw��1�oo��n(Ӭ�O�̧G%b�!�j�8Ve]Y#�u5�����4|�-��?�O?���~?����Xo�������9��5��4�se��PO&��'O6�ww�tC�EI����en�u.��E�6`�qh����%�
"b:џ��T�L�1���/������k:5��ƙ@_Bw��H�B��=]~�E����Ӹ�J1�!�V��Iٜ؂+��&EUs�*LgP,���с=Y������������X�SY}��M�:�[����h4����|��G|����z��%$�Qm�M�ea�8b:�Y�ؤ�z���p0�&�U�������Y]���O��6��^��2@�1��#M��$0�3����8�Nx��7ih�7��i�u�8k�i���Jz��m[f�>�W��'������石��Z �^S��)O܉�H�	��=�ٲ�����C�Z&��G�~�d�MJ�%I�D-��{�l:�`o��G��y�W�^Ŕ�<`�����ȓ�S.]�`4rԓ=?���_���~y[s�-�C�%�W�t��<3��9��������;��F%X����Z+m}H���N����.��?$�DU��5��
�;<ԓ�GgL�O�N']Ex���͔�B�ޙDY8o��`o'�EM�F��)����������{��x���6�g�4�Y�+^�Au�?�X�f:�Bw~����Ε,*��\5�ӻ�.c ��ͨ�MTeA�a�k3[ �n�h1��jn��'h�H�"m8Z��s0> ��ԶB4g&��ۯ��x�YM���qHS7<Y�I����b����|��|̅��
/�=+z�X7�	��x��g^�+��j��j��N�)B�FA���$�B�	�������8Wa� }��'|��O_A��W|�O������'�Z;M��ǅ�ֶ�ș�Z[��¬��{{����Ҷ-�ᐶ^tԀ�E2��dڏu���L)�jV�cz.Ѫ�aT.����򓟸�
�oO��FkL/������Ǒ�2a��K�U�K~~�ӑ�ib��e��{�M�����E�tMy�:��X��I˞ږ���o��	>}9@QW� tm���Cd\O�I����0EC��)���eg�)��Ɏ�H��~�ij?~̯~�+�<���o���ϙ�p�|���"b�1B
D��:�������<�~cZv������LC�s�ٳ�,9���f�����p������MӐb���t�Q�&�B�S�*�����=�pv�W�Q&��_��S��Tw]�[���L����s��}.l^"Y�`<e<��g}�2kÒ����gw�.O��gz�K�BU�C!�x(�l;�}�8RPB���f��?�*�)�1������|����~���� _?%�O�O���Q�@�DA\�X!Ɩz6CS��䰻�)6� :E�DDsG�f8c(J�T�^hSM2UK݌��W��!�m���o)6�EI]7�Pж��aN���C��RN���C��b��ռ�p��f#]�UL!��8����:5�K�gP�XbP�5X1(	M>��IH*X7@����b�Q$Ke�0����̅����-޷�~9g�j����]�[�����O���c����is1/��: 5�b�y�W���fw����[�1ѵ6�V�vXɪ��Ŀ[8[��u2����a8����G?����_���'vs�q��?Y�5����?qI�'�A1����4m9>8ܘL&.�,�D@��<�I��Y���`�8�f�����#�N��T%�:��lc*���*$����3���s�U	A��$Uc�(�|��E'�~��S����C6t�Wg.����8�V)�k(V�#���2�޿��8�qٖ��U���~���k��o<��_���t��*�k���f�	|M�cB}H�v�<��d<g�g988 FK1(1����;��1���~������|����6t�-��Ɩ'O�p0>���#O[�3���-W`��6�:�_7��V����>١r�������JLk:��k#�@��hB�p�ϸ�	dm`)�!Ea�}"�-e�!J[�����c\�&ԖH��!Q�1��Q�QڀȄ䧐��I!���1Xk��@���)`�Hg:]O�k���r�)�Hf�А��Y���2�m��bPr��JT!h�$���qW!D�`�v�#崣��H��F���lJHu��i�mZ�R�1B�&Q�HDf��WLYfB�<�u�o�o�{q���,@U�o���b����͆�JW@�L�����lC��l�}�I��M1`�ҕG*�mC@	����{9�|>F��F�9��YK���/:0I�d޶-V���H1��L�;|\��*^���>�;vrn�[D��Q/�$Ĵ�
{�IBJ~�!�XSUv�&L��OJ�X����~b~�㟙���gG�1������V:w�R�ܞ��c���z�Q U���Q�g͠���Y��#y1*2\��qQ�x�X�Or����j�uSծ�KlLq���`/�n���x��,�O�����L�V�q�&��5	�N�-�XTɓ�Ƣ�U$w��<,�Эf��)�m����Z�F��lfk
<-�Xc+�t<�Z�����%�P��w	�RT�v���e���>`K
r�1M>8�*�4�1�3p��{�7f�ʈd*� 53��Sf������}�n����1J���8��!�<��~���se�*1���ȣf�)I)�6?15����ȕ�
�1ⳬ����;�[��bp��J�9Mn�RPtm':i�j��-.�rv>y^U���sʪB"[uV�i�c��l>/H!Rh��~�ՙD$c��su\�P���s�6B؁�C�����>R~}вh��#��0L'm78J�Ďc�1� ��@Y�m�����'H.͏_ �ݙ���EJ����`�J����:��^��t�-�o�!Q0���S����k�':�N׵/1�<g�.���UC*����I�4�'����˔U�82��{D��k�Gl($�^#��WgX�Ou��EP
F4��巏�Pu��q.%%H�R�5�[�H����I6W E�y���\���������7)X�)�|DT�K�f�W�RJk�&R��f���؋&��0���J[��+��O�n�?�ѧf��j�w�����S4w���n���'���R��*�K�1�}%�������U����d�1�r������A�ˆ�>t��������?�Ʈ~iI=Vk1)��)ϯ��Q��L��11)��@���Jj�0Ŗ�%v������gc��U:F�0&%!�u1�d����u�?Z��7�JB��}CU�y���(�������EvN�/?�wqH)Q75�{{f��q�����n�V�����
!t��ɼ[ċb�ZK+������r�끗�*(�"��B�٪Fcw� gW����i�$���V��G���O��8�~��U��*Q�:H�Y�;c�F�����Kg�.�5��O�wf���p��7>�[Ě�K׸������>������I���6�E��m��(T��!������]Cz�0v�XhQUuRu�Y[M7�f6�!�)��d.��^/Y�u������t���y��������^}ߢ8[!�z�=
'�ݚD��d���_�+8�]��Z�I	��]X�8�w�����S�5M�d� ̭WV,Z,I�-W�j��X��+2@��<~����]BH81E�1j��@����!/^dss�A���0�����$3Σ`����O�ǐ-d�h:��B3k��$�:*5��XYM���2�8
0^%�8�����*��i:���y�&��͓�����1W8ۈ��v���%�d�q��GEQ�����ч����_�6������U����pq:������z�O,l<']��'��>dk�謽��dR��ު�쟪�7+����!��)�Z�j�4�l4�N7Ƈ�E�4Y*�V���ŽesW,��E$��I�(DT�ALix���'v^��-�3rlI�HL;/�:s,"9����]��RM�QJY���֗���A��>�X�*@c-�a�h4��+���kvvv8<<̀�Ȃ���t��]ڼ��o��[W/�6Ќ's�O��B_|.�Vy�� ��++)!��*�3�v��\�����A�eA�:(8��������5����?����o��=��~˯;��N0�����4�+��ê*�Y�F�U�O�[8�/[�M�?+Fͧi���TվrՌ~��?��ʁ���w����?���>*q���?�,������U�+_i�FwyjL3S����b+�?J��7��w<�[냑Sgdm0l�1ƇP6���Y]�O��y�^�ڟ�Si�_Ac3Ţi^@�C$��%q8+��ί6���<^y�Iӷ���$�I&�K"&i�����`��;͕&b�nA��� ��a}m@QX��Q9�og��<a{{�}���x)2UE����K��" (Y���>�r���'�������VX �$Yk��9�|ik��׮r�������Ã��2O�+����N��F�����lQ#�pe��>-���E!ar��ף�>�W˓�d�NJ/����4�uX>!�k�$�F�Q��j0��?��sM�j ��i�Q.���p�P����Ц;X�����׳bˇR�n����z�%���vZb\�&4��8w����}W�vW�ߨ��ٌ4���������
6S9*�5�~���v�b�Δ�rMqV\ҤҴͰ���tR�,S�[u���h���~��@5%$t ��@Hڦ�T��^��|����:rxo�Pp	�6%HJ�uH�9ӷ�^~*ɵ�BF0�!"�͌���\���/_b8(�~��Ç�~��z4����6j}��%�b�K������ds�kX'�f-��v��E��5��iU��$B����pĥU��qx����cU�'��42��v���i裐��T����x��_�3�|���q����*Nf�~w��� �o&�������災��qϩ*Ei��i"EQu�z�m�Uj�Z_ۜj�֕E+FRR5)�.!}��	�}��~
��Y��^/�֤Cm�P��G�!<����ڎ��ҍ�{ab�nĢ�k6��B5ҡ	0�n��6v͖���?֔>H�ه�UAGU5�UY�\TM�o�Q;�mx�}�ڦi�v\���(���&^������R�c�6DB�F�[��y�o_�	�ŵ$d+�؈:U5"G�ď퍗{���;��#����"]C��K|��;���[\��"����Gܿw����K��}ȕq1k�b��(��P5(��Xc}4��'���=e�`/[6��y{�{*ٹ�ϻ ��    IDATH��Z�%���鄃�]���2�N�L�T�����Aa��i�Y�TL6}�k��1��'ѐ�0Y�>\���4}��e:���E �U|���y�5^���_�G�"��Ѣ��N�X��DFeYVj��� )�PT�ںn�1�^5����$�=I�`�Rnc���ZQ�E����jU�q:L��D�Vn�GFt+Z�D��tr	�+Q규wkɷ�c���n8W���Z] �@<���:F?�L��I����t:z��|�nKO����{��.lI���FB�4��U�I��1\��~��� �-��i��(`�}�$�dR�6�/T8Q�Ē<��1	���)Pcx��5޻}�wo\g4������#�>}�o)��ި�8�̲)����F��P��������YSO���:#Y��-��N0I��b%kg(��Id��4������H52'}+i�#^ F�bD���J�W�e3ꤽ�����w��v_���y�&��b�{�%215�Y@U(܀�pHJ	��_��E��u���5]S����R�B1�)�!�Ԋ�Z7j̄H� �u4^ ���v]�#����)m�&�a��� �c5O.���cw��/��2��\��-��\���E�����B!M�b�{�F�|��?8g��MqЗ�>.�X^�d6E�PD�pe]W N_��wOP�ڳ��FM�2\[����*�!�W�)x��w������7x��U���޽�l?~ȓ�;��I$�eF,���	[qEE�F4m�(,�{�ׯ18,���|��_�gUU1�L(\E�b!��RG�+��	�ʕ+8������W0�1�\~�׃,�
  ���������r��Q�ٓ�2 㤮"�������<�D�wg�A�	���q����}6�s{���,Kʮ7o۶�I�vZ���/�����糂ھ���kW�ɯ4��L심YN)冚��Wg���.8"٨:!�h�����{ՠ2h�j*�"8gP�2�Xi�/$R���V�zM�Ψ �
�*;�ͫ�%O�����P8�jJ���0�8��l4kf.���s���ׇ������;�eM{	UW���}v�(�K�l&�>��\>)�}0���ӟ&�����[gb�Jk5U���%f	��Iz�>�~�㪪HbH�-iC.�غ|���y�;�x��UF�����}u�P�5�]�_�N��j�blژH�FL�ŋ�q�m޽q�A阌�9�ߧm�DB��ш+���u�(�BdPX��u6FCJ� �L'�L�����1Z��	�t���fiۅ,�Wo��t�LC߲k828<<<����8�}.sx�at1$r�a5��<��E�)x�Z�h��(E�*I��S����El0֥���8��AEDEcD�dj��q��)]D-�4u�&��!�!�*xoC�4�r�Ƌ�u�S�����Q�1j�Qb�x�cw�)��MN^���`�ٲ��ֺR���}A���XN�������!t�Ƹ\�Q�z�&|�޹q���!m[s��W|��_���}f���a�D���*�������n��wo��kW0ֳ�󘇏�3����1FhB^iI���GX_��z�*�/_f}mH�3&��1��H)��p��/��=8�Mq�r��z�
����8~9zV�(���k:�3�Fͼ���~ Ů7�t�|�ShE0�řO��[�5bR�)*�@JEU4�I�Ģ�k�.�;n?+��EPє��dU�A0�{������p�{s��߿��Y?rQe�;���\��N�<ޘ8�{\�+���M!/uu'����5Ε`
\5��[7���l]y��2LǇܻ�_���ܹ�%��!)eX���	\��� SW�+��pĻ�����=�~������{<����l�%kQ��I�jD�ź���$�j�ƥ�Wٺt�����a:�g6��O����g�!���P2�v�v�V�|��Y��x��h5e�c	�'�E�ӋS���X>7G��]�����}�CU�G�f�y�Ҩq��������+FZ�5	�$�FAS���hcD-�I��,7�l2(J��������rG�|���ӂ�ש��x���`�1�<C���!�կ����gf����RKnM�]A�Iz���j��h�(�؂ \X����~�ÿɥ�ˠOy�����_����<y�M���j:���C����9�5��ܾ͋�����ryk��-���<|����'���]���U@=V�`�)sJ��`\6v����>�Oi�Iw#�\XqV���g��i]l�	����c�oE,�{��ih�����ى�П�k��+�����-ֆ���;Q)�B94�1�5�1-��`:�*kr_�Ō�<�Dke��]���5�B�V{����^���sm���?�J�"��:1�
�&����˷4���5��j"�eT2(S<]�]P�P)%bR\Yq��M��}��Zcw��|��o��/Ν;w2���PK7X/��ՕZ
g��իW�y�&W�^�,�z����~�ٴ��˒f1|���N1�`��Rĕ��FC������d�����b<U��G��J�JZOڞ��{�}ľ��w��}�D�D���g.����)�+ˍ?��`��YW~�Z�1�3,)ET��Z;�Є�[P��<.�`qe,�Cմ� ����~r��<�e��ke�Ln�YΔeiLW�e�I"�ꕽ�y|��L9�*
ߚ^4yU#�X�dR����EE��X���L&5o��ۿ�����Ν/i��c�
��v���T��\�����n�s��tL&���=�7��>�i
k�{h�%F%���Մ�܈��%�]�εk�p�Ѷ-�Ovx�����pn�g}	Ë�Az��㟷�J*I����������W���X��	�������%D�Y���[��3K�v���8A4�l.߿��x_�C π���U�a�x���}Z�3���{��&vټ�M����9 ��+\��a��j�M����� �㍎3��Y�)C���J�b$:�Ϟ�c�cK(˒<@�d2k�������9�?`4d����5�Ic�����[ܺu��W�������Gܹs��;Oh��Ҭe[c(�2�#�V��x�"��~�o_�(
�Y��M�Ǵ~�R!� A^A�9���j�3}ov8����=��nguss,����e�y�=�Nd?�U�K_%{�u���=���m����Z���.���4����z�ε�0Z�I�}ǹ�,�g>��8F���8W`l�ֈ�5�	��@��_�}�'���8��#$I�Ĩ��Q�ѨI��6a)vb��� u�>��B_i+ �S���&�<^��?=���m��wvA�J*¬��D�x������O̚@U��쀠`�a�q��[ܺ�[�(�I�<����|�)���S���`��QC�<X�X���Q)����*�X_�k�����/�՝<�W�]E�Y���t���a՟�ϼͫa��������S+��x8I3 s�`ur6s.u�������wr��<.��f���7�_s���v��'E�w�y��O!=+������7�#�d��ǴB_���cN2��O��%F�U���ZO�~������IX�-tL�v�M���Ο��Y��;�,�Wڑc=p�}��N<[��2>q'�I H�\?��7��z�K��)��x�^�[#��-6�礟S�T}V���f�g�2���Y�>�E�j��"�=�G�`>/�Zͯ����[f,!�ު�tm}��f��pΥ)����v�j��ε
ߢ����'PL���|���*�����}>|ȝ;w�]��SU�gQ+F��p=�L�ommq������u�666�L&|��W���?�w[!���tt� 1yF�7o���ߦ�*���r��]?~L]��f�\�����߆X�p�N���~�-H��y��=��޾�����ZyrtBx,�|F%���O��߅.^��~���=��n�>���Ua����[|�c��҆E�/��U����M��,�_g^�Ǖ��� �ˎ_�;�qΉsN�u��uZ�����������[_����O��G�7-F�VEE� ��r	�Y�}JJX^]�̩�+����}�n��'hBU��!e9�m2X[[���?�>|�ׯ_�ãG������/x��q���ɫ��Bm�^�o0�aL�h��͛7y��ﰹ��d2a{{��>������4�{�@U��6�"s�on���e���Y�d����X�L~�3kF{;������߱[��a�Dt��Iz��d����㣽��n҂e�N�!��g[�*�}��l���&A@���nU㉠�E�A���Y>Þ/�c�AO���~�o�?�	�y��q�Ӥb��eP'K��J�w��V����cL""�\a��1Xg���f�{.���;��g��ŵ<�%��Ր�GE����VTU5_i�1���
�f�F��v����8\�(�� ����&����G��7or��E��}>��s~��_�t{c�����$h�%З'����Wʲ��[����y��m6/l�t���`�����Oa��sߞ3}G��ۣ�^g9r���:�*�B��(_o������:H�Dn�t\ ��|�G�:"$zI�2"�������j&e��벤g��N���.tvϜ�%����2sܛY��+ow��'�Ó~}�ذ��>I>Б���2��S�����e_G,�w1;h�􄉱��9S:�ֈ�^ӌ���'�g?��Y���7(��������kn�E?�b"V���?���aޝ�B�Az��:?I�H�m�1�N�!�u�oB���o������;����ŋ�D?~ȧ�����/�~�F�*���ӗ�ж3���ck�"7n�`mm�m۲���xrH-�r�u��r츕ٷ-���8��g�o��W��93��m�Ukw,_kk^��<y�Ư׳��������g{����ѕ���u/<�f̋�N��%3��9�*��%��J���LO��=��;���<����q,�i�(���Eq��x����z��獛}���U+�Vމ�Κ5��5�����1gouߠ8[�ݢH	lJ�`,�d��|c)g�5�{�s8W�W�ٳσ�&3��^}���dp8��p.�ԂZ�p��%nݺŇ~ȕ+[���y��W_|ɝ/����!�� �ퟮs��|��������?��}�֥M���p�����rZ��x���m��M���c������� �\����X���z��"�x��BT>?h��$w�:��L�gX�W�<���3�)�F3S*Bf�̢�d���*�3�ǧ�O�J>(DMWh����J�m5�������~��p�5�Gu\���ī`�����^��ιcu½��/ɋN�2~��3}=��3} )%��.2�IuՕ�!�J_���/�E�g�g��
<�oz�	���|�.�n]c�4��5������@�����v,�8.���F�2/�7�t���\��1��Xm����p8dww��0�����f|����E~����e4z����~��U�i;cP�q��{\ڼ��H�6̚)��!�������]�dQ��%z֖ q\��i�h!�|��&n��8��K�z���>ޕ8���h�:�x��ǂ�[-�XT�0��^?�>��`�?~!(Q��,���*^���4��o�xn�����vL�1�9��@&溾�LW���@/<���7��5͋Ɏ�� p�ƋX��|?�}��3��2�{��nk��lB��Ĉ1QL(4�ʵ�����y��ę@�A�ɉU�D��"�d^�:)y�������u����z�*�������s�c]�]��bTK"֔T�u�p8��W��x�ob��`Pq��%޺z��]�^7��)�lK)�A��U��>�����_��_��w��`�x����';s��=�r���f?��f��:)��0b���q���Y��*qV& =�͸�N�xFW��
0����XT0ϋ����Ed�0'k��V6јȋ
5�=��~�Ȍkϼ��~��ǅ��9��90[a:�/�u;�wʉ�(����۷E�`0�,K'���Vq�)��y|�����q�����q��Ό�`�w7�ɈD1N[�$C`��r���{�3��ٺVZ��aJi�.���b4�{����2��_��'�bLs˓����yY�x��������ܾ}�����r��=�nr�)��*��[J4	Q!E!%�A�d˖6,,)$��|N�>W�Un�|(s5�&8����o�q�-�~���i3f����Y�|��OO�SwmI��~��
,L�v,*b�-r{&���������q����o�3��ߥ���TP�2�ޓ�Q̯�����:4�4E���}�]Q�l�_N8=/b5D�6ʲ�G)�:k��Y_��o[�FՀ�t�`�(
�4�(*Tc>>���!$R
�k��q����٬�mg��e*Wa
�GЀE���!N�X"�f�w�p8�mj��2�͘M'�豦�үB҅!oǀ�����%y��My��!׮]����?����u=/2��)%B�\K/g�?N�������|G�r�`+��:NwgN�W�uW��>�s���x߫�a�x�[. 9��{�Ngh�c�e�|!�е��DD�X+)E�օpoc��9%�-��i�fE�d���f)�&�Z�^D�r��Z���d�����۷y��	?����������"�7BϞ�Ч�\'@�H�!��	I��l�Rpue��?�ՔMl$�ّdH�`PJC���q��gO�9��#Ƙ���G��ٌ�F��⌥��X�4&�&R���!	�*�2�̍�B@K��A%a�+[QC�<p
T�+�d�`l�MCUX���/Ė���p��0&���P�:B:�.6_��A�#�,_(܀�j���W.1(]�ڰ����A�A�.P*)�"��#	V�,q�0k[|��x����d����F����t�C��p�2><d��C=~�ݯ�dg{�Է�R!�|��m|���{�_�N&=z4����<�GZ��k��}��܆�cY��鋗^^.k{����}�_�g
U�I�y���)�0)xx��b�ř@_;D��+*��;�a^b��%-m�.tƂu­���C�Ww�`{�EQ�������Kz�QG���&�������RV�M��W�^��$_Z�,n�UJߚRW������ɘ��`I+=<�������>m,�����6`lg���5�ѐ���J:�)�Õ�XT@c"��E�G�쀌���8ہD7}$�u1�� ���	!q��8�`I�����pPRV����䐃�]��'��|2�F�g�k��$��Z�ZT#I-��z�mnݾ��k7ؼ����pP�֕���iIE��4�.��*)F��Ě�l�C �@���T�ӥEQ ���T�m���Y=�+L�Ϧ�v�{�����d�`�z��2�t���O�}o_�������m�+,q?n�)��q�8
��_)��#����8fO櫲���{��y��V阽��E�ͳSG?��N1%IIŘ�ˈ��%�ŤP�&��s��-��߆�Od�׿;
�fC�j�>���8z#/?�t���{�q��E�������]����={�c��j5PUU�t���3�58�0z=N��L���oy�fm.�*������{�r]�4j�V��|ٳ~�q��I7hb0�@�E�ePٺ|�w�y�˗/�\���81����`'S8J�8�N��� &#*W`
Ga,�C��R�v�
+�Pƹ�bĊ �RXK+Î�2�W��1=ܣ�M��_�����3�ݽK�	c!)�W2鉭>������r��������K[����&
+�X'x���dM砪OU/�[[�����l>ى0�-X����Sȩ�r�ƈ��d��c���K&�CrEr���ު/�s㸔~ߝ'��q�ެ}����.zP�0��;��X�[8��yR�g��C�`(�b�Y�:����~	��Ԉ"��1u���Ι��<�aq&���j�J2h���Y���S�g���C�����6k������K���� �� �o�DoΜ+��Nu�    IDAT�~b�t��-ȀO��u�EG�gW뫃Mh b���ƐR�Z?C̳��E����:�~�cy5�� Y# �5�߼�����������¹��Y��0�m��ӿL�SЅ�����K;k�5�����93h�d=!BH�	p�r����e!(-)��+���3(+�z����������}m�C�؁"A�d0����[|������w�JH��{8��$c;p'���c{V=����wk��T!%Hm���&��,WR^�AE]�L��y�����$i�$�C�D9�����f����n�Xb�z x2pXf񀕖��鷾S�r���o~�����х²Fo����Ξ����>�{��)�Ŭ��󽐀F���ak��oz�q&��xo̚؂�u����E���X˫�eEJ���ڵklooc���*��)�锭�-��X�#�1��~�%!�Y0��������7e.� �~G!���I��D�8︐o�g�=]��9��2�e�Rg�c$a�8Z�;�}��?��ܼ�n7��-��&�0����w��$���~k���|Uf��ɶ�vђ@�#��2<7m5�� �QNhX ������dXMK�\�$�Q�U���s�#{������dVeuߪY�d�s�9'N���X�[���8KflB�C���`|~��?�c`D�T��1h��D��=](BU�)(	�u�%t*΂�w��!?��S�%�m�	�)�yۥګ��H�J�Đ�3�pr�>�l���ږu۰Y]��\a����)gGt];�],}uCUUx�ǂ��9�v�ۢ>�FXT3�K�,��ߴ�]~�fu���
���r�{��sr�.��,�Ec�Z?��9;A�D�u�İo�>j7E�4}��4# ���_�M��LGz���ϟ��y��@��T�=�g���@	U�mۑF0 ��V�?_��-h.3c7WWw����V����f٭z������3�EU�AS�2H�w���)��r��M��?���DY����/�3�2��j��A�&T���ВĚ�B?p�y�ܸD�0ҧ��$���B��Z��ڍ�����Ik,V�3]�wb4U6��ng��{c<<�*j���ܽ�wN��\A"���-�͆�=.�(�|��E�DM��.Z��'��ɳb�(xLヨg隖���eg�m�����ق��i�5!�d.2�g,Y�ʲ�,K�ީq81D��V�k�t<���6�e��X� i~Eeuu�'?�	?��_��ZQ��|�l��ݎ�n����iƍ�9��n���u��U��m�^������Ȭ��v�_^�ێ�m *�|ƃ{�y��#���������yA�X��HBL�(ߐ�t��~}�����4U6�߾����noo���2ӻS�~�y�c��(�1��nԑ�78���c�}�ѽŶ֎Ǹ�M��a-�1Fڪ�1�M|��wX��"�ҧm�g��ɒ����cdou��m�VUE�e4MCUU��.(˒�(���O�{�xæ�{���E��l0i;���'nR�7'�(�L��5�C&tB7��!!�q��Ǩʻ}ᛲkW��*�O�Ӭ��eYZP#�UΫ/y��%O�>e�^�c�\2����}H�գm{�lY����� �����v;b�cZ��:��I�SeWoi�5yn������?�Xi|U�!&�k���"�6�>R����(m�u���:ʲ�w��}��������3�2�*s\~��n7��*�2�����2qз��Ib��뢌,yq��8kH�����sN~�GGG\�ڂ��W��w> ���/��/~jbS�g�T�s(0�w����c���&�L	y�����l6c6���y�!�}�@fzb��X?$|� �Z�EQppp���"���%��_�6Қ�y����V�������l��e��l	a�FC�T25Q1� VL�$�F�l�/`��-�G�)��]��0��-�ŌˋWj2�db��M为��u�!�	��O�tp*�Hw}9�n���L�J�l�ح5�e�Պ�jQ	]�fĘ�֊�%=��a�!xBƔ��"D��;����m}�)&:����Q0�Md�k���#\�!MS�n9\츸�S������_��/{��"��Ξ�}�����ꞣ���@`l>0q��آm��)�G�T���l6�N
\~���.}tD��8>��3���M���"˩��3���9��T��Ѭb�
��c;f�3*>%^�	���Liw�t9���)���eH�t���D�03<�4#ֽ~�D�JG��iS��P���q��`�6��yEYΨ�/Y�~L\,���[�q��_=�i���-���R�O�D�Z��a$ �� _�ٚ�l��k�ը�ٗi޺%o΀|�N��e���Ƿ����so�o���ӣ#%`���"��c6��X,F	��븼��*��?ZyVrx�����NNNn|��޳�J����w��%����9�l���]N�RP�Y,c����^�FJ��������wI�<~��jQI[�.}ݬ"y��k�B�M��g����r)�ٷ�n��8o��jL��AEzd얛�@��G�T�s[�
��~������&�@��B��zE��HfY����nǫW�X.��y�l6c�^��hQ�F���cS�\G�M�pvvƿ�w?���ǜ���L�=�����{P%���C��I�)B47
5RAG��>��&3��:T��A#V�lh;���6^�z�j�����+�&vTT%�_C/^���v}���c�5j��	�?�,�ą��"��}e{��9���1�Rц���3d����?��l>�mClH�ж5�F��L�k.�/�;�[Q4M3r��|�]
-`�皻�K?�u�z������r9��<y2�?�٢k;88�v W+ EQpxxH�D�躖���1�$�4�ۮ�3G�ٔq(���2�q!Fc��1Ħ���:Z��ڭ�^��a���(��g�F�og �j��5F	�O�e9�U��O�Q����URu]ߨ��3l����T���1��u�͆�,_C ~{���m�
���c��gϞ��9�g/�!�����0�`��`"Q+�S����I�����91��V.z�`%K��%����h�c h���l�k:�`L�EQ7��5�5L:��b68}�MDd�V��7u����U����:ɹ��z$���d��63dY���1��y��[C^��yI���w��c7:|o�K}�����wk��g����T|xn�i����'�s�{�= qT_�z5�iV���@~ѿ�$u�!�%���,�'��!z�vsE�����bD�{�k3�&�6�=m���4eI�ACZo�Z�ױi�X҅���,{�Ӗ�Dxxg����wYU��tƒ��T���״&ݻwoD��-���!b���$�O�~�������n���n�b����HJ���M���iޯ��?�E��g�=�vOhۖ��3�;2�rK���x��W�&IC"���\z1�yyC[��܌�3�#��[�!���,�r��$�#�8g�rK���}�j�BO`z��a7���C~*=-f��,�XT)-�.!�m��5�> ���b�YƤkS�{����ϖ,���������3N_��nT�� Lc�o��eY�/{��%��1�Hc��4h��x��c:��N�8���j��}ey�>�I_�m��)]�m?�R�u�޽���GD1�gC�)5dYJ/�!��������� d����%��:x���	�W�{�5��j).
���������;��[o�r�N�68c��g���*1�[�H�~�P�sb�cg����־#���AlBp}M�ZK�&h}�\���V+b��e9:�������Y}gߜ����AJ��u�j��$��#f�� &B�l�:IKB��Dl/�# mDTq��ӴhD��p�<�)
�ҡ}1I�4|v�&�@�j|��f�Q�@mWՃ����yۊ���;������]�α\���}�sBӱ^�i뚮kGt�,Kf�YB�eH�����Pۓ�]�s���#�=zD�~��r~�v�����g-7Rh���;{�y�o
{LQc%���v���?��?#��f��
�<����ؓyz��ƨ���\B�CHE^�md��b���{�r�d>���l��j��wt�����	t���JK�F|װ�l��ի�^���jeڶ�U�1�"���ߴ�s��|�~�w7\]�����H�zo��ŝqR>>~��<~���7�?~<��?��c�裏n��<~������e�gv��a�QA�(j��w;ޑs.q�4N�p�T4L�餚���Ӷ�f<M�0\�N߳\.������|�ޚ��#Qގ�M�9Mͼs��y�"���b��w-�'�*��Q�ۤYB���GQ�HJ��Mڐy��?y~�PcZ�1��ƪ����rpp���)�|��NO	�ë%F����!t�\��؃[����::����\ڷa�{c��n����,���p��14�=��9UUqpp���!��h������5l�[�O��y���;w���rvv����&��%�J�e@�Ҽq߬S�M۔�2�wH�W�/�N��S�n�������l���Ÿ~ܤ8��=}(�@��8��n�_Z�25cb$�@�<p}?lgm�������W�5��2c9_pz�k3|�QgK���n|������y��v>�}�C�1���U]7��fS���Yu���V�������ݝ�鳏?���9|��G�������g������Ţ��=~�<~�8�'�m���u�e�������Ν;���ivQ��|����޽��������#��n��_�f�7���Ǯ[�_��?��r=�1�g���V�7��3�ϯ���.OO�Ν;������?��G������ӷ[�c�\z��0�p��(��Sq�����S��w���$N�3gpʦQ��Ѿ��n��e��'��T�,#�k=-#Bf�3�Y��2�K���]AL�!����	��Ȋg,wf��CUU l�k6�Mӌ�l6�ZKUU|�;����1��?�)?��QB�/m$�X��M\f!f�eNQdI�y�0i��.������9g�HS
9fdƎ�5�Z��1�W.c��sxx���]�,��
1���eM۶l6..V\^^��/�dl6>������y�=e1c�7c �x}f�Q�o�������`{�k���A�|>�9w#m;Eꦭ�Pձ�p<�1]ō�6#�eΠ}�zP'X����u�n�����ݎYYrtr¼�(r�s�*X.�{�=�+	��{���Xجa�3�����m�H�F��2�vm;8n��X�t�ģ��Є�;u�y��k��(�J��y/��$���h�����;��]8(�͂�My8߬����Y�i��E�m�����D���_�W�a��޺��f;��J8V;�{U����q	pڿn>��O���v'�[���Ƥ)�F����ٳ5����QY�f������w�Т�,�F �ЃI�]��֫PF]Gs$&�F#b�.�5�|�
�nr5}�J�h�0qI�,�vW����m��*)v;�c�U�pJ���C�u����#��>����sk��ιxvv�
�z�O:�R��h4�)�u�:��ؠw�����N^�IL��i�����������,˘�f8�n�o�F��}�q�\������kS�}P��T�������(����w��x��W�%˃��,�ˤ���|NUU��\�s~~�f�D�w�y��}�s��~�{��s>�O���3��Qr��V�^Ƈ4S�%���0:g_E��m68}��5���!��Jz�\Qi[�v[���Rf�jVb���9稪*��B��[�&İ$#xO�D�6�B�Gc���.��!�?�O��ǜ�]�HUUt݊B���f����&��w�E6� E1��5M3�]��ƈ���m[��-����|>MӼ6��E#���=X�4]�y�(�����G���{������#>|HY�����](�G�wPv��H�O�I4��Ū+=�_Ί��6Կ=��e�Uӡ�klB�ľ7�ZQ5ǉL�ƴ�Ĉq�U���(�5;1�V�.��F3+f'��,l4���D$X$8�A��UT�ݖ���HMl���hT5A4�5�v���fp�ҸZb�]yﵫ�0""b�����I�D]�z�g��%���:2o�ع�Bv���D�Js�p�!*�TH�M���K�F��f����fM�	Ar

�QP0N�yI�1I���9�s��U9���LͽJ�.S��Nb���Zڶ�9��J����=[����a������M��VN��ё�"��,DAMT�FUׇ݃ߵG��S?"y�KS$�3?�|��fLqu�'�_��5��?o�*+��kz��?��M��(�N�(o� d?�<=����FUӁo��E�ݝ�7���s~[��mc��ɞ�����3�#|	�-�kgJ(X_]1�9��9!��6\]mȲb��ʲ��|���]NNN��"��("4!�-(燨ɩ�m�qx�./_>��/���w����٫Wx�R��m��&�,�y�j�Z�?}�_1lR	Ŋ�3�!@����ޝy�Swqԥ�+����|�٤Pe�������]ץ���yY�u���"��(�˄��,G�py�e�kX�.���e�Г��o���Ֆ���@3Ќ��gcZm�b����.r$�<U�����%v���u�r?/g���̩��N�����N�������~�/׎H�n�%[��Z��x�#�y����� ��M��#%$�4���f@���������~����srr�Ç9::��@w:{y��t����Z�+�]�|���a��h�]�_^#���
11���FL��J��0b�11m���9uY�5Q�!Hf]$�Iʈ��� ���!�����3E�r�X���8��:&ؠѢ*�˽�]�dY^;��!�1b��ykmK:�`�M�mTTՅ]�cn6������	��jUc����D��ֹ����NUQQ�>�����i%5� jhDE�u��X[���:5]1�N���}�e;��Řh1�d�S���Ҫ��l��Ζ&���Wͮ�;;<�7�9�!�+3��u�e6k�j���������~�O�������5�o�@*Q��bT@}*ݠ@�I���.^ב���i����y�/B���T�'nH�"���Q�e��iï7u���OӖ"B��d8[�1�O#�%x� �A�\ˮlYg;|��
�g��W��@W̉\9Ǹ�g�Ny��W���6qآoA������1Ό±�9�.	['_������&��S�N�I��E$z��M�qxxȼ�06m�����n����kܮN�]V���'-Mo�\*r���W�����9����?����S�#��+���!�v����e�t*{P`��o�1Ӵ�4 ����o��:�y���c�n���!������ܽw��?>����|�ᇦm��ߋ/x��)/^�`�ZѶ-�k	a�:ٔ�*�$���ը��V�\�;s�Q�80*��x�J&J@�1�Vq QP��W�8���b��F���	^�rk�WBhQ��q	Ռ��n2K-֥�c�P�N�O��K���Y��5	~�C׷�T���}x}���m���Ö��*
EC$X�(�^�k0�͊�	A����2'�K���D4�BX7Ω�A�s�Q%FED""Qc4.˼F1�]�fm����La��f��k��<8yZh�c�w��3��umϲ,<���{�����������_��g"��r���rG�d�"�D���5Q}��N�0=�yD��?V}��u��7'ؾ�"���h�n*��6$e�#����۾Y���ĩ���O�����"_�l���X��"6-� �q��vӢq��6-�GK�,�f��>v��nP"B9�Q7���1����?pvz�v�P��w���� ��*(�GJ���ucRAI�:d�^$i����$ۍZZ�a���޽�F�e��f�P�%�K�'b�46k�@���X��Ҷ����s�뚑�:�?;�ɧ��{v|t��W�\^\�Q�?A����_���w����3��uh�o�L���4�3�7E�޴���!�5�J�4���;�-��?�GG�ѹL���cUU�m}V�Q��    IDATo��V+�?�ӧO9==e��"Q)\��D������Ԣ���Q;���+T��!*ɿC1Fz=M��Bc����з����j�9q�I�� ��	>`Ħn;�K뗵L�HU���1�nHE�&����±�w�J��1zBPp���*j�WY � E��@�j��XL�R�V��=�c��>!�"XcG�NH���HL���t����� �Gt����::�l�n��� b�GI7
C�X�GU$�2(�f�2���B���lV!F3�nU�s���ф��E�$�>{�������)����ݭ:r���uf�UjF�"����D��V�.���}K�µ0�t�o���C���������L�!��&���^�����42��T[K���,*P��E �@e��l������A#����@���#n1#���y�:�Ѿ3�Ř��9�S^�x���Wt��g�o8��̐;��\oi6M�v[|r�l����ٵ!�lL����}�o��9�s||�G?�pQQ�9���ټ�	�7+�%	}A�DM�I��ƞ�\Q�I��NB�EQ��S��� �H`����=��v[z�� �n�՛�~���?�toJ����Lm��,"c����>��C�����w��l��IloBTӶ����l����'=�a�z�S�����;���l"�b��R1�1���1!
1$�I�������1d�%�=�!ɤ%~VD�`\r$UQ�e�z�'��R�y�6��x]U%�y��\U�_�3Ϡ��0��u)#��<;�����۶��U�����`��%.'�]ZK��I��7�6�X,��QK�$�.l/�o��q�#���)H�#�Y�3 bDpVȲM�o��\���.#�G�;��NRp��Q�U���,���{Z�Z#�m���A�U��E�a��hu���+˟֮�������ӧ�[:}���j)")�TS�a��`H�nzw���+��_r��|����x����}�E��@D�O�����ЫwHߛ9��ocS����׶m����kG'�<z�}��>�Ō���2�ȋ
QC|�ֲ���5D�����8�XɈ�ӵ����W/h}ǃ{w��J���\UE�#�~_ץ��r��pq~I]��e�s��"�or�n8Q!@�c���~�*����C���!�������O?O)h���;��T9]w[ʲ�����y�3����w?`u���┋�s�֗d�cy0g�I���t��;{g_bӖk��=;Ӟ�S�ox̀N����5d���b>���������k��k�����t�3޷�Xʲd���牎�bS�D�P��mi�Ժ�w͘�v�Z4ڸyTET1�H�;�H�{G��A��W��(�'��[*����c�b��J:N�-�mI-!&D��_�D�5t����~t�Āok����it&�Q��?ט�®k'1F�bUN�<!v�TK�54J�:U�ś���8:"VA=�D�+0N� #DA%�XR����)�� X�I�u$��78k��tmHWbr��]K�Y֑4�u�6uhR�wl-bL:�oO��ɜ��Ǯ�|��I�y!�*bT����w�l�\)aU��s��r+�om�:@��,�����)G=���kT�!�����GNÄ3��k��-������<��S6���/�h�vTr��6]0~�׿������q�&Du���E�&�����8>L���ܻ�٬�{��1�.ru����n���1� ��$+`�`l���F�6Pf����.M�c^��+��^^D�4��l`躖�z�sx<EiF��� ��oZ�n��z����b�����<x���lF]�\\\pyy�u2rc$(h ��������'M��b�ɝ��*��O?��?������uMYe,����e�o䝳�m������q��=�{�f!���k��s��y2���s�ݻ�ݻw��Ί�ԫ�+��ù$�rqq������zX���Eǖ�0r�� �wF�	����9푿069� ����8�O��Ǻ����9@��e�	!v�~�!�{��:���@�u����@Q��5�O�FDL�H�9Bp=Zx���'�SJYBķ���x�1gm��r+1�H��!���&�`�D� ���1��D18��N!`A#���TH� "�9m����}.K��	tɡU�RA��)���c
:�4u��E���֊��k%7^M���/L���Q�u�uB�l[U���?��?2�J��_FUU,���TS����熿���q����.�}��#��Y$��$�v�t{��	��y�o����z��u�:1s���brH��~���y�	�w���T��\�k74�������@���=����X�E�`1�ٻι\����3�N_a�b�z�d�Źl,�0���dGׅ~&�/��u���c����}��Im	����n���+v�K|h0ɲ�5}Sy��Al��+˄V��Md����%WW�\\�%�2"w��a6/��¤#���;�~g�m�Uy�c6��Z��9���,�>}�ڸ��}�ћ~k�(�N���u�f��x�����L4�>C!�o78�]�h!/��~D�i4�E���2K)M��b{dӆ�'�T�Oȓ:))c!��	�A=��	�2V1�@��X0=�-e"ҹB��H܀��y�-�әQ=F!�*�IB �"!^#i`ȝE5��U�I�T$�J������Q^��Ū>C�������t�1H���}��ͮ{���5�K�֌���ǙaL��#y��|O�a_Je��з���H��ش��kE�����Jg��$D/Y���mp�ʖ!/Y�����:��<���5�}OU4�$���]#}İ����_w��& �O�������ސ�"���*��_��6ٴ
z��~]�0��ZF���@��lVr||ܣUk�f�fs�z����ݶy^bm�t�&E�=�Y�!:��i��*�(E&, v����ӗϙ�f=R��;c��'�f.Oܕ��ӵ1��L�;֙����q���+�>U�����������2�I��Jfe����w��O�h��̲Z�X.�TU�ԑe�횧Ϟpyy�'�|�j���'�����(R�|6+�w���:}?�9���X���~��Mg:�c�Z�l6��ݻ<z��}��k��ӷ>Ӡ�,˱��v�5+<x@��R������ *�H�ԗ� U%�^���`�s%#CA��%�D�����ñ�Z))%���(�Ӎ�؀s}#��WC���Dm����������'��W���i�����G�ff�Q ����%R�Qz~�D�I{p������{��m�
Ltt�?ǌ]� �$���\WYw��Y���E<��8��~��)�Z3:s��er�D`�X }�i�����?�8��EY�g�o�.���&��eծ(�:������ό��Y?�����ٟ�ٟ�.���J�ʕ�]�ԵA]Gɦ�r"��Ut1pqq��ppp����3��,�����7#�c����!�?��2�h�%�6�T�c:B�ݘ�S"���5�]�I�_�1=���M%ZTu�쫪��t� :�~��qkR���Q�9�W+�(����%.�8>>�Y5�C�����wPu�OgO�c�h�1Ĥ>ف.M~c0�al�n� �:�EL�䁮k�tI�uc:��̲↰��F��K�Ǜ��B=���BE1Z�S�i�bT8樷��`��eX�"��C���6,fs�Y���9�����k./ϰ�p�H���}�v[lY�-mӄ?<ZR��M����sv�WW���윧/�\�J��|A{��/W4u��Q�a;�qii�qBQt�c(ˊ]�b߀$O�����_{H�"��T�)�2U�)�Iʹ�'�4`5"�������5��N����]���ã9���E�'F!XG;���?��c|�l�5E�H᫳s��/ħ?��������n��a��k2�:�.8t;d�
�{�*�n:Z�Ĭ�n���G�*@�$D�د�W��:O3o�m���_.���Ͽ]�T�U��w��?����:Y;��h8;����o�#%��-&z�A�T2:brB�W[	X"&v=��}�,K���m��|��/^��,��ΑYG�8C�
�،�_����U��bA����1<z��|N�u���s������%���ylϰk����(�T�d�X���Z���+}���T��y�5[�U��!
��d����wԈo"�$U��H�q"i�	�����z7�A�92w���t��9�~����+f�*Q2d�&��@�Ћ��y��ډ)Ö�*� �'t�=��������_ЈnS�u�	�"�Nh��8�n�g�q��0M��7,Ĩ��WW����t7)*!]{Rv�ZK�K��&b5�������|kC��4�3b�X�����U�y��*ۧ�=��;���=�����r+���͑9�sng�e��7�?4ָ���bq������ܫr||�n��'?�	>('''��?��Ç|�;�[��ЦJ����f��>8'�A%r-r�����O�"���(�V+f����5a̶mS˜/5C��uUUq|rw��l��5�1de��b4�yvcQ��&UI6)�����4"�FޚI�J}z��K	��!��}&�]��6p=��sT���O�<��'ed�&n��Ʊ�D�e4�TM�׹a���cK2#��>����3^�xE�4x�l�B��������w�4���PM��Wu�SN����N��i����yV�>��qyy�RB:�$F�r>C$����~AA7�o;DW��PsN�v�<u�i�@��fGizD3"�6�a~��:���s���v|g�1%����D*�jO��:ƧGTԠ�;���Ħ=�m�)��(s��Q�A�y�ٰ�6��f��?E����}$i���ck�A��իWq��=���z̦
�r,�����M��6���qy�bWo��u�����9�>*1�^��5�RV�Y�o�njb���Y�(1�� kՈ�h�k��"j�ب�ֈ�tm�����.�� &b�11F%��Qɫ�'�1VĊ��%&�;l/�"Q�=�$�b�%&R,�ԀŰk�t�%�kɭ%K���m�c��#�!�M�PDERn]DDQcDȋ�!�:��V�h�ѐ�� ����$I���DMH�pbF���(z�F|[L����<ύB�#UQ�n6��ƽ:�l�3���Xt��^��f�uu�Ύ�Pxa�絬Vw�����>4��#w�]��Z,we�>]mοqy1__m���#r�.�͖O>���G~�_�:��[��~�������w����z�n�A�������c�!����u�{|ұy휦��s�7����c888������a���8�
�?R�;�IE>F�(�E���`$�/gE_u1.E$�7�dLS�)e.JP����װ6�C.+�6�kS
q$`kPZ���_��NSb7y	�>��zр�I2���'O>���Ã%��"��K<���#���c�ݎ���� J�yֻ���J"�����iȳ�!Jd�l�ϒ�rQlv�XU�/*��6�!�(��Sn�v���oB��3�����QV�jFQ$��#��A�+m͚t]c��a��u��imC�4dE��{��]��A^���Y{6��*q�G*�TO]�~�_�x�u��&�� �o�}�:1�����}u���LE{�A�����{1��!D%(X�1�r�9�����;	���ϟ��:!���z�}��^r#��0�^��NM�ӛ��m[��i��w�����GwX,c����fKV�D�]s�WWk�THB��qآ����A��^�Q5Zkk���ͮ �!Q�Zc%`�F#.�P�J�(i�S�F�� �ص�c0BT�h�E�ɜD��x�,��Q5	8%WL�Iu&����h��|L� �C�EoQE���C�ƣbS����'jp��bTo���Mu&����D5Q�(*&`Ԩ���^�DT����A%�:qV%D4L�����de~EP�ZŪQk�$�K^[P0Q��D�"����Z�}�pyV�l�n�?���ؼ��mk/W]4��ZSΗ/c>mB7��;5���ms�`S>}��r�f��ɬ)K[:g�u}L��ϖ������<���'���<����������~���<�麎��'�>�����z���:���uz��N�x����nJo��m�ޘ��}����X,������v��7:H{�Q�+�-�_�xfՒ�,8>>����fC�J拜��M��(g乣���,+0&�cL�Ve(�W�}$���e��-ƪ����[���q�y�˗�	[;�\��'H��p�wbBHZR���4u��O��η��-֤��(�4�6�����Ǯ�����$�@S�l�[ !�yVpxxؿޓg���<{���nGY���'�P䡿�~AE�1-L�˷�o߯!�r��}�/ƈW?��%)�Sf�;ܻw��|�^I{y�Q��a�|��{]��g4�ѣ1`p�����C�1�Vk�.׈���)���>�W��x���_�o�&"��篻��M��N���J����zA���j̐�����$g/�ɆÚ��ڶc)ˊ�G����|�;����=�����m9??�B��m^s��Nݾ�K����hc��Q�%�Yjƺ^�YoJ\Vp��{#��g�~���Ϲ�����紭��k|�gs�>�2#sE��U��,�X۱\΂�U\�bи���^Y�M����T7�1DDB�k'-5�0FZ�N{�R�bD��a��B�@�E�5�5�1#�%CU����Pi���AU� q�gD�H�C0�#ј$ *�l>����(��b�H!ΡN�LP�1�^@}J��֤�a4J��	"*B��Q�`� N�1"bzb���+`D,j��DL�1F��g8��N,N}aqI�P%KM݂�(Ɗ:�PE��'bTd���fWKS7��U��Qe���(��b��˳�6��6N�%&����]G��p���s�x������ӟ}2����Kg������~���{�71��gO������}�v�e�M�^�I����h�D�b5L~��Z�q��d������ hŵlF{�s粛|���A����������ײ�J����s��E��Lf��UE�%�n $j`�p0���x$�dO�T4�&6jJ���p�$��b���.����ͽ�t��`�}�7^4� �ɬ\���⶧�ͷ��ַn0M��@)�T->b��������.ZB�hm�T��+}�) A��(���ֈ�dD1ZU
4Zg,�e,��-m;�,�<xt��>��O�;Z�9��mFw~�2�G�a�m��Dƌ�(�x\���Ÿu�![Qr�y�eͣ����{�wSd1J�6��~���8����+{W�&��O�N��2V꬧!(|!����>x:��u��ǆ�A�0�%� xK�v�g̦�NC0jz!P"�$G*�	��{0���+��'�8<�zL�^ 2�E��2�H���4�?�'�'p�B�X,z��k�������Z��{~�q/<���v@��٘[�������+/�ҍk�l�@5�'�Gg.���m�6ı�8E"=?�u%��r���w�]i��<�gP�Q|����G�q����Ѡ�!u��>����k����1� ��D+��4@�_�&�"w&�m[;em3v��V���^�_B�6�(�\���>�Wo��V�g���Yk��+Wx�߿_ ܾ}[������Z��U�:(YԕX�ЎGE8���s�oo/���$(��tz �U5Q(
?j�6.di��ɲ�g��"`!4!�U"���ZP�NL�MJ��B�.Z' M�S*(+$�SBy��RBz/�tN� B�
1�/�`��2�XQ���B�P�F���gI0��R���)8�C0ʃBH!\�W�hB�Z��,=ai�.�M����BdƁ�o}pn[y�-�HJ���/��?F΅�y��;����_�B(u�>n��_�u��ڰ�f����2�����)^=?<���ի�x���������ʫׯ�����{�QU����5��M��Y,�H\�|�B�8�Z5U���J�I&� ��K���F�ןdu�P;-)D�o����J�_�.��9�~�u^}� �و�i��ڢ�sF����Ƶ����m��^"�    IDAT� *�B$8�d�s1��\ܬk��1�B�ՆJ�h]P/�@�#���ݽFg����c)�M�W��HV7"�
8p�&GQd���5��ªRQ5��%�t����X�4zW�Z+�Zi,	�zpF)�(��Ҷ�Q&��<�E{~&�1L�'N��1O�6@w���Ma���ה�EN%B�vL!X�*^�Qn��,�~�C}��(F�gG�h�����
�c��,/O'�����i�,�9���g)W��{��	����OJy������Y���_�����$?X�V�����X����]<FE�	R��d��ǝW�ɛ��;ܼv����іs�Y�q�ڵ�/n��|�����K�,˲��:ڄ��f\�������S/k���9|t�|�$7��tʍ�n�IE��`c�U��ٔ�h«�ޡm]�&����> Bt�t1>��/*����k�e+�:w���xY��g�TgR7�1b�_+���?�hƍ�r����]k�r~|,D��HQ��9���^-��΋�B�\V2m��cW�4���u�T"����)��-N1*8畲2H��W6x)�t��ޏ��FFI�*��J
�#��ҝ�,BK��I�U7¤V��A��R���U\�Q¨�DV�m��C��؂���5%����F{-D� ����+�Xu�C���<���uP�U��B@�&_��̜��if'�X��ű��+j�r��F�Vu�װƸ�mE���kN�3�PB0��6-c����@cãr��>��A�X,�G#����{�'2����2�̨�^��7�1�����?�?�z��M������X�i������,�������'Ҷm ̲��֯G9��'��l�N�?�#ȡد�'R1*��)�.�g�c4s����]��|>g<�!��F�1�;�ؖ���oq��mv�v{Ep�c�"���f��%8h��
�k-���UJe��q!2B"���{WnrkQ������}C��U���K��1[�X����ȁ�9�q�t�WcGJ	JS�%mk�.���A�<� (�̠���-��($BE��YI��
���Oi�$��e�/�VI�j��l^�x\��ƛ�� b͐�Q;�6���5�[�R��_i%vV�(YAH�X���ɶ!+[[[�y��������5��3�v<YW f�f�R�8E!E�۶e>��|ޯ-Ҝ�m��o�6�Vr�خSB��I���u�D��	�0���d��yԾl,m3����5����������F�&h�|���	����h�����b:����#|�}���)�{�"�3E1��O�� �m9:=c2��d@*���q1fk:cgo��x���uՀִHB�≕�A(���U�B��Y��A��Ω��_����:�3�te�e5,��$xӜ��4AklfDH)d�/��Zj���Ef����J���@��"ӍkE�&���a<��E��)R/3��v��j��Y�V���@.sh��Ω��ZZ�h\���-弆�	x��m0~�۶�ң��^kC�
�@�(*x�ڊ�P�IW*�t-���!����I�*���RZ��.SN���{�H���VZ�s�\ȫ��:hmCM.�R�;���0˰�b������ ȂZ[8�E봒N�����a��c�\:)�h�H��U���L_׳Ҷ���I���K��;�^{|�Xܽ{��J��G?�Q>�N3�n�\���rY���ٱ?��l�_�1j*W��_��)u����X.z~C�XQ�2M�E;;;��k^~�����<��h��4��HD��r	��y=O^��}�(Ek��ҥQ�aX#�h�h4ekk�K	[��QV�%�Ķ2EV d�m%M6�s,DId~;�]k,��Ź��ֱ-�{6u���"���qaPz���
�٬O5A_�f��ջ�HY��6�d:�!�+c:�,��ei0&��Ľ���n)�U��K��B�|�]4Yu��-&K�K�Sb	���*�?3�S��9pP�L�	����Ǉs#�>���n��,��0�8�r���n�x����Ŀ�d�w�L�� e���-n߾�1�b�c�X�����x�J� �{�(@/d)힎x���_Ş���W���"�08M�(놲�T����P�e���y�[,��|�f��b�7��f$=�yyv���H)���fgg�=�1>�ivv�z��ml��-�A�0�c<˘Lf��cw���-������z�eEU5̗͠i���ŕ���|o�ʃb�5���ն�vP�� ��(U���i�?��?�������cl�?��?6;wv�ݻ��ܽ{W�+�<�n������ �O���uM.��\	������t��6���ݻ]�6'�����׹�=���x�Aw�#���Wu��c����R�E&��t\�Z��w�����?.r9j��s����3ᔒ8ȥ�Rz�XN�B��.ŸiJi�N6۪�B�|ڢʕ��m_��p�p2/r�Î��K9�b\
�j4
EY�J� ��U= ��)�쁗R�u�hfM>�TB7e��,ggJim�k������'����ޘ�F����\iSN5��,F�O����������m;���G//���GcJ�+H�ܽ{W�����d0�a���r^~����'ׯ�����>0����-�,ʒ�|�U���M�s�jٮyI)
�@댋�9R(��":aܺ�{04䞥��1�:���0z5|]zm���E%���W1���Sc)�u��L%�Uu��/*&�	{{{��N�\�}/Ҷ-{y��,;���`�i���S��PJvi�mO;;�loo��k�`kg�E9G����ׯ_痿��ZK����o������X���mۧL��y��F�NJ�X�1������$:�$���R��D>����,K�g�ϳL�#B�8_��5e:����`��6F�mF��W=؊Q�؆-I!%�d=�������4ϴ����*Z����I��4Q�l8��s��z�F1.2Dp|���<|������_�¨JȾ��t�s�\L��0�IU-���f:�0�a>?gR�}1E����%���B�P&R���ӚϺ~�⡽��l����阓cz�t�P�uEX�������G9]������ �4���.:��PUι^�nx^J���";U��c�ұ��k0�B)�K����4���E�W%R����svr�������7پ��:fY�F�ؼ��>����`r4�a�����O�1,�U_����˪{�h\�ل��bL�:>��I�����ߋ� BD�����j:۲U]����Z�N-����]�����O�n�S�4h{�O��O�B�w���@�v/ ��Y�ON3�d��u����������~��B�&=��m��+���������w�>����+ ~�_��O�I,����],�)�O~�Ez�}��������L:�&*��O��Z�{>�������&��𘦶\,TU��m�;⻖Q�$6�o��|�����kO�mگ�n����Sۜ��	C��&l�� V��H�nBNN����ϱ6�����9:�(��l���6�ٌ�h��2�R,�K�m�P�5��ؑAJ�Σ��ry�w-R�.*�N"�lo]�ڵk(ex3�,�"���׫v������o$��1%�V��R��r�����Bj�#:N��zK]5ض霅�P;nd�g�e<)�(���K׹ru�,����d���y�8���
NRt,�x��k��;<ݵ�a��%i�]8R����cGGG�����7��|��(-E?߅ E�dq.���>(|�B���_�E>��
]�Pֹ��]�>ϲ�R����v��5�N��Y����&��4PI�V���Ǯ
�E�s��+_�KW@V)��CXkeY�<���ixmdX�nױ��#�Jc1���,��w6��9#��"���T�1|>}��a�.!��j���%:�v����\\,8?��kAz]��Z�������y�|hl0:ڹ ���8/���_�n�W�~@�W�$!�B����֜R���-F���%�V���1.+���B5ֲ\V]��AL�@�GLR4 .�q�{��;�Х�:5!e�_�S ��FA��{��D�u2�����_l��%1�+�)���,�Ƈ�׋q���R6Q|��M��Fi��He]!����a���=�HK�u�tE�E�G)cd*h���J��/�~��n���x�=ί���s�]��@��$>�F	���qH�2����<x�����s� :��ὥi,�q�2B!�Qp��0N��0��(2ʺ�:��b�G/,� ��qL�&�(��]�$��b�/����>��s`�s!m:m�2?�`~~A]V�F�ј�Hk�u՝k�c�Z�4-��<Q�5˺BJ:0+x�]����Ż�������_w��߄םM������5m��@��C��/�����#|��E)Z���!��Tb6F�2��z:~���] 9 p��o�RA�R��i�
! ���T��s4�C�6ri۶����~s�F��OT����'���:3��BPwm���$�_�٬�gi[��%U�62��U:����J��"�`�Rʠ��� ��r#+����}/g/�͸�A�*쎔z�;ޮ.�j�[��L+#�m+�Hmc����������lş��DN�[�l����I�䋤��퐿�*��b��~���փ�T��-;u]����5��x��A�Q�͒�ىo��ki����L_���x!�"D�hO��-	�&��E����c��l_٢�� VU�_�H<�L���bY ��u�x}%��9QH�-����Z"�Ƈ��A'�#�z�T���-R	��<2�6EⳮsN���{R��E->(�Δn��v��0ґ����&�֚<���۷oRU�pzzJ�ƴ���IN�2nܸ�h4�������DG��� ���N�`�S�C:F����Ն@-X�C���k���4��}l}:�����f�Kkݧ8S����UJQ5yV :�<:F���YA��H�P]z�B�tp��^?��2��>��-���N�B�H-�
�����n.|X�9���t,�
�aT3=��J�h��&�7=��)%]���|�|�<�i�lL\o�~J�a#0M=uE,8�b����� �B�B �]�7��_�	��F�Aߏ~����VB���k�Dx�\��M��=��r_�QMc�VBi���	��������,k�]!GU�4sXq�I�O���G�@�u���@_��z�=/�K��fD#mr)�eQ~"�z�`a�֚z (�x۠��f~qF]��#9wTh�rk�t���"dL��`l�-K�����N��Y����ՂE9�n+���X-�k8���_F�R�\�0W�ù(vj�AI�:���}l�����،<�jg��w9*ʾ��Z�����=v�jI���`��ԇX�m��M;���"I�Em �}#���j���#¡K��o ������tʝ[���%�lo��3�Q#D�f��7n�e�>���������n��R�i^��|���xM�9̗��Cp�����ۜ�B�\nC��#
<��k�ް7y_������ZO�bb�4�d�QD�*��*���يk����f�A/���E��#GXE�D !Bt���*��!F�Et&����ԋ<��t�����Ɇ�z��4�ctUB,KiݢXU�6�W�~Ew��ή�����>:G���7"/�pa�r��Ʌ_�WԞ����?V��Z�L�Z_�PI�}�loX/F���!h��Bʖ�jp6V<�e�b�`�\R՝j�`���gll��GEV�6A��ؐ��;������nO�����i#}����HBFmom��=��~d�8P�Kc����bR�T� c�B�ض�#��n,ZOb@Į�6�M`Q-�M��W�%ی��Q���۟됬�eYWuk�wR+��նu(�P�'ޢ�D�碦_��v�z�.��c�g�/5tH6������ �����(� 6\�s���d?�g����lm��ٙ"$�&S�� XJ�u[��LF�Q��� o-Ai:l�G�DQ��:ܠsI�δQ��˾�%�>R�v��xX���@k�^d��=+z��J`��[�	!8??,0��%�p;	��<��{�W^����N�^k&�(g"%k�����A���`�\������w���i�}���k���/t�͡�v��m*lS�J��º��u�2'{�;j��s3���M��a�_j����>��|�9�v�AV?��c��N1B���]1�s�{'D����E&�pA��?Uw��w����ϔ���i���K/�d\��ڦ�i�ۡ�oi����1�MdB(B`�����CU�,�Kʲ�i�ޫ��L<y<��|��RR$.ti�4!C���K��~ÈFz���5ӂ7��t7��K3D�	�u�5Z!B����M�S��6ѳ�]�^A���m� d�<�9��6t���bU�`p�%�g(=[Z���]����^>�^k����09L������%�R ��?�w��9�[���g��l�z���k+����Jhvw�0�ls~�����z�!���b��m�@a�jx�C`ӟS�u�����'�c�|So�����
@�llϩ���{7�1���w��Z�CL��h����G�M���	e��;��u�����Zں�>?g2ʘ��\\��qqq�����8��iKU̻��ܹs��7o2�N{�����J�����G�qxx�GĆ��i6��Y�q��-^�u���h۶�qxx�9L�OgyT�t!T�'&�-��*�����ʕ+loψ}������dru�9��!��߿߯ǩ:XJ�Gע|�YbZ4�@�,MS�45F\���՘N���4�W�<U�.պN�H�~e�������}�C)���	K��&�)rYe�g7�v��<���  ����',�K)�T!��)������e���!{&����Ea��B�.��M����ŭ��!d.�Y�ڶM�P5�Wl�4\\\pvv�"��{z<���a�b�e�͎+/h)�>L�$]�M�aU`\��?p��TBpx�ҴqS2]�!.Tݿ������RH���xD�F����Wd��Z���ֶ����9εa�F��Ǐ���REj:ס7/���d����{\��G9��]�"���=����X�� ���Ǳ�(&�|�\�r�G���s||�Ėa�'�6��#+_�ml�������z����*��}��� EH2u�I��X�y��}�1����y5M#[ư\�,�
�$����(u^r�:����=><�(88�k�"�D���d���-i����|�����7�d{{���^$�/�ܿ�w�}�>����}���Z���lM�N������?����e���>�������=g3����&r�V�h�x<�ڵkloﲻ{��l�U[�uG*��6!B�Fݤ��L�yN�\a�!�/Yn4-�֦}�Ź����=�6#�J���x=7��%o���=���E�}��5]���22����{��%�u��g�Dk[��D�TȂ�)�wNxB�k�����X��'?�r{H_ۯ͞�*���ۚ��Bη��(������C�~{g�:[�mB�z�y�E����t���#����JM��Y�e����u֥Z��fк���NF�U�}3B2�`]����)�#P*0�Bȼ����2��N@+R{-O� H�!r�\@���Œ�j�"�;�"�׫���=��#�ж+1X����N��B#��X�AZpb��;hs��\ń	�Y�-1£q=A^"A��;!��b��"����Ł�ӿ��T�W@ ױSIE�5����,>�m^�l^st���6�RKPc��tdN2��A��l���.g瞳������;�!M�rxx�T�(�4
)A����Z�l�2�Rh$���8�dΣZK)v���b
�G��GT�#\3c>o�׊2LX�#=N7�� L�h�/tu���ʣĂ�{���������	/����#>�茪�bUMۖ]1��i���S�F���A�!	,|p�#>��N��ͮI�1ʵ0Q�i�αl�����Z�Lf����    IDAT�r=XQ�l�����a[a/.x��}�|��5|��G=�mK\��"$�o�^�oα����(�>�����!o����(]����t�W9e�
��h��#�2
�y�o3����_��w�-����_B�d�s�&к@���AP7'y6��+���0�����{�G���y��QL����¤�c����O��ã{d��)Y��i�[��	�;Zo1�m|0\�im9)+�|IiA�]\�chj�4[ܣ�-�y�#���-M�E�����O??���9���x K���K�+32���~YU���HtW���Q���Zl� dF��ف�ʠZZ	��u�[]�%��p_J�Q�d2YE���W��L�3�`�$؊Q����Z���m��]�gu�PE+����'~���5��v���O~�g���F���e�������m4��mS�m���qV�\ۚ�r1�"!hk�H�ZY������t��S}2��i���<~��'m:�M��I\�gِ?L$sί���+%k �@7��--"��I��e�����ަ���8Kq\���pzz���9��"�r�_�o�w�R�[[[L&ڶ���,VC�RA�-u]�eLM��]pzz
�����t� �F�u9�1)
����0jZ���c�2X�%��R�bDEM[u�4��9??���ggg�(t@
�)�e>,UU�ӟ����^��������^A$���\�� �Eɣ�c�j%>�9�6��Y��_�6]���1J����*I)�N�YN]�#���>���G9���|�"�D�n[�f������(i�9�~x�G�c�Y$��UJ!t�����9;;�W_����=�����ƭ[�\����"�
�����ߡiJ��k���=���lW*�aEt����޵\�ٍ�����&�=�;WؙL�'/���n8<<���}���p���b�������et��O�~}�1��dC�4����&��2��g�&�h���v~}�4������<?�=��lD�N!��cc@�	)����Tq�w�{�m[?Q�|��ھR�D��o��y�P���������>����y�|欕)%�8��2��I�uC�Y�n��?ib=m�]69�mN���0��<�g|��6�7\��0!�m�I�V����1i��X�f�{��sH��z�*����P'��x�ˈ$!�?����}�������I�t�fdQ�,�cggg�����>GG'�Ŝb�Q6U�Df��޺��JF��8M�s0�C+�4�}C�<��P�������9:9������R��ô/ҵ�ƴ�!����Q/K�}��-B���� ��K�p�tk2��o}�;�nvU����s��d{{�k׮E���'g�<x���t!�����4K �����~CmMc�n�m�_ҡ,�`6�f<���t8�y�`������cL�۶�J1.F\ݺ��{�Ř��өb�&�)gg�|Y#��
.��he@)������|�{�����s��U�Q1c
�� I11�~U#��(m����()P�T� ��,�|��'����f3�2(�3ݽwx�o�Z��Ԓ�(�m�g�~�/~��}�q}.ж5�iim���E	I��]˦S�i��� ��5�`����mF�6�线4X9KB���)�����Cǉ}���?�������f1x!;�2!@�y��|�h۶m�.���eO���y�PJ��u���������U�^�u%�i���n�z���3�c�/��I���?)�&�����z�M�˵�ަ'�����=�t�B�����$�O�(wQu'j��V��<�#}�i�=�}�-��C���^�@���0��w����"�z�m�`%��$�?����i��T�����:23��.��f�j���"��j�Nx���6�4��9�E.��0�B�0�I-τ�Zj�.]�,U=_E<dlٖ��>D����j��E9?���u���3<x�Ғ�r���)�����C�b��7�z�:��'a�)�Z+��7\��4�֪`���,�x��Ke�{�TdZ�n������W��/x��88���&G�8}kɌbR����~HӾʕ+c�f��x�W��u��ѽO8�#@�LNn��X/OGl�v���m^z�6W�^�+�r���m\g�D
M�%���w�޴-6x~��_�����xo�ʐ	�ف�����T�9!������l^���j�NNN��_�����?e����;/R,�����p�F�n�t��)�r�7#zC����a�m���y���ק��/�qY�am����sx���ވ.
!�A�����|�*���w��]N�|m_�.}?��G�,)G�r��<7�}k�"ǅ<X[�U�ؾ��m���n5���+B?	����`6'³#}���gġm
i�k�T���&hn�����3-v�h�"�i��7�҂��qn7���'�����)�KH�ٞL���6̛�
��TfB�{���I�%�E��/��<�p��������)Zo���KKY��pq���I<�'�g�<Rx$�Jx�z�s-UY"���Ѻ�T���G����nh��E=%#J�����cQ�?:��.b��!k���2s�_֑̿����������Q*� ]��1�!p��M�wv����{N��D]6�i�g��xo���Z�@��-e���K-�����Dmȶn�R�<��9?��ˇ�>�v���@l��#׆"74����|�U��aRL1f��Uv��"��X+^�4��A*�����[������Ɉl�̜����G�89����n��׸ze�"����o��Q���S>�A�Hap>�Enȵ��Nb�*99:`<���������-���}�O�	�Qt�5�9��E=���#x�Qp�Y%����˂CG/9C'p3�;�5x�|��eA�V�Li�Rq�w\�ZO�򑻙���� �y�k2!��!��}�i/..��/���E��I�>U���fu!��.>��=��R8�2k]�"y�A�tΒw�Ti,�G�6A�����'�U/� ���'�Uz���n�06m<��u6\L�����M��t��ӳi�s��9���@��@����0��#i�)J�e#cG�t�����soC�{��(��>V޸q�o������IPU�Vv������#���� �7�.(��3��F
��l@k�eTu��);�>�(f��k�LJ2[
��)�@����)���T��ց�vR���˷��-B���lmm1G�7�N�������D�.wP�|2f�6l��MkЗݒ�L]V�4�b�����hIP� =���P�������2����Lg�Qڠ�F�����G\�q�7��m�����;c���9����+�������!3���)o~�[ 3�v�dň�_�;�1ϸ��<��n�Jl"���r*DY�kj+�]KSW�u	�#e�ZVZ�L�ZK�mc�8HB����ȠR���:��63J	lmfAV�T�&ْ��Pӵi�����w��a���;��瓢|�<BH����(*� ���]q` ��T��/���9B_�W�}o��vѶ���#��*����Rd��s�;'���d˪�5��R Ն��:�2�7�'EF�'z��ϻ�Ƕy<���_Ԟ�"H^�Uc��_������{~<GÁ7�?6��.Z����>k[��b�m�l'�b[��}J$�U7����k�x2����h���Oxh[�/N��BjW��˯F}�N,7����CzK[/pv̸�L'�MC�ZH�-}A��(+ٽ}qԧd�

.~^��l_A/�,D'D��\�޴iꔢ+�G��ҭ[\�~�����6lmm��=������C>��s>��3���d��R�9PisY�����:g�!1�&�b�O?/|_к�-�Z��#��<S4�pX�"���.�������}˻��:Y�ڠ��z�:CX����;�����?�6W�_�0����'���|��y����G|��4U���n��c<�p���L�S��#ڟ����#��drL$�E���6Ff�%3D'��%���K�H|yD�*�S�&�s�ZE����/��G�9��^�o0��Q�˲O_��n�����@��>����JC:A��د7�!RI%ʵNz��!���l�/tB_�W�}Y�����N��`~h��V��Xj�#B|P���\\�b������ڶ�ҽr����j��\О����_�'�Ӣ|O����MI�.W `��6mC�Q1�.=��=�mr�.��<��y�n�U%o�e���]B`�D��޵έ]��jrP�g�EH0&c:����KU׼���\0�M�_q��+\�v���=��������R�������'L��'��e�s��N�?BG1��zįA�nu\2F���ƬG�AU!�`�V��D�SO��0�DG��U�����:�m�N�r||�2v����ˊ�j(�&�d�b>_P�j��������zd��q����i�T��� |C���%A*>�
���e	�cr���	�~~���9�o]#�69٨��k�|L�O�fʝW��|����=����:��䀏?|�w��w��3*&h3bY9��'ܫlӐ��ֈQ1�(
2}��ͽ�?���1AI��8��5��:���#eҿ��a��a{�T��[,bˌ�}�m)�k׶4my���;�w��	\]f鵛���Vlϲ��!)36�	�9�.=�'�כ�/t��Y�"���
�۶�vޣ��(��J[�6~���EQ!�L��[���·+�h!����9+ j=���Ӯ����p�X�QC	V��4d����~�EC`�xp J�~�%��m��S
�o�tC�LmZz,�K�RvZ������g%��������A|�^j�7Y#D�3��z~IU-㢗�]�2��\�w��	��A�:��$���J�`mۢ�^S�-��@�����W=#��燭�ڶ[ػ��m�RQ��...PJQ��r�7t�x.�%�~�m	��V��ӽI"�1��y�.p�����Y���"j��lw�t�ŽO>�O>A�N�΅���P=??G�t:f�5鮅Z��q�	��xa"N��x��8,�HU�����Ti�e87攎�R3M��ܼy�s��atN���%�~�9�Ucx��7�&����,%�ɬ�F�e�d4��D�X��|K�$�eS�yF��(�춉�i��j�B0Oh��O�E�G�G�@�#�K���$�P�5����!(�b��3&�)��S׎�7n�ƛ�ag�!X�Q�x�d��?x��G��#S#�o�1�L�8?��'q��o�v�I�G 0o*�]��믿�{}���D�ڶ��]d`-!8��h�=�}w���"G"��e�
i����MS�ܬҠ1z[\>+/i���Ul��/��D�e����f�Wi]��Eֆ�9Yz<��9}�����&�iHQH�6�M)�Z��dY���jq���G!��#2���Z�P���t~t�:�����dk�oZ�Fk-�.r���͵{�ry� ʇ@�C|6+�`5���L�o剈u�1�w����O�e��
�o�f�ox�c�*웑���!��;'�I�����t���]��\��7a�]�a�Lj����5Z�l=��&�����w5nW�b� �Ĳc����)3��lo���͛�<ċ�h�sx���~�s�O�;����3�A�B�9 ���)걊\���}!���9o�c�2�qcy���|�7n��g��͛�w���	�n޼ɭ[/���e�zf��8L�{�c�E�%s��n1Ҵrpc$�XI- \��'b�G�G��cB
�A�h�L��B�T��#
d"V�m�x��u�'̗%J��b���t̍�7�y���%! e�ֵ?!�'bJ�!E�:e�+� +P4�Ц5<i�^���q6�6���(CN�e���|2��S��c��K��9��|:.�c$4�5�S}p��,)�����5���F�CX�Z�f&��[o�~�<������������n<��&�����Jd�û�!a�����ZOUU}��չ��5�N�%���$�#V�ڢ�eY/߰\./%s@�	�6%W��>zR�q�zuB���wi߫W���&ppp�sm����s�{�1�F�~[�oӫ^'���6E)ʴj����m܊���;�N��൑��X�9Ej�dy���yUrpp@Ӷ��#~�o�u,l0
k�Rj�2��������+��L&���7�:����<v�H}WS�7i"<{ %෪��w�v/�T�l�M���C...��f\�~���6U���_���l6coo����_�����-�n_����'8��m���XW�����.8l��@J���:"j�I�q��k �Z#�J�,� �֝p�H�Q2�輏�`	�fgg��~�����1_�� i��m$�h��h�k׮��K�����-��(�8օҤH1D �틄�,�c  �߀��W�MD���k_�Ս��_��۳��X~���\]�gR6�POs�7���a��y�e��!(�cr
c���Z��8F��b�M�I!*˼Tm^
{��6��N�Aߵk�dQUҵm!
�mx	P�����&?�%W���ٝ�{>FD�SD&3IV�J]��%Ah@���� �hh)�J�6h!h���$�����Ph4��"����$YIfdL>��fv��{���##��,�ٴ����xG��|�;�q V�ng!�Ty:���V�N�q��"lӃW7f��.rڽ��`a�:)���ӿE�J�Q��?W�����
�?L*C��:\-����͛7{q�rqqA]����_���~���?�n�d|�M�}
���c�o=S7�j���-���s
�v'�!��u�,�8::��F���E�ц���s�3���py��~�9M�k�&�US�i������_��_SE^Q�K��of,����k ���/q*~0��������y��	�����w�]�x�.W��]Ĺ���d�ܦ4UU�u}��1-�َ����c��U��� @�F�"%�^���_�d>M�l��1Ɓz���FR@5����X�'-x�iRpt|���w��Z�� � %vr�|FQ8#����Vc7�`�Ez��S���i=�Ȁ�+=�A�b�%����1FT�L�!����^sJ@<��!�X�D�jp>���N?g��+�p�Z6|��w?wwN���S�]��]���e�����bY�V�1"��k!�x�
���8F���Gu���_��?*l��������hT��2�!�6u��M3�<��@�Ո=���y㺛lhV=M+�P�e�NlW��:-�ˀ��Ŵ@�Ĥ��tLA�"��f���i�X��B_��w۟籧��1�ئ�v [y��Z���)��P�+�v��x!�~�>7};�=���+l���4-��~��|�;X���ϸl\f(\IY��tng�o��&�~�9��4MC���0����t����4�����U����.1�7`��϶��}�����l�S9�T���Y��uC���s~�ӟ1+g�G��b�prr£G���@2f��WdW�]�}zs*ȏ=K6ݗ�N��-�q��&*��v+���5�w�}�b�%���fB*�Qk32���ɞ�e��4g��rA] $�؂���Ѕҹ��_�X�f�%�!�%�;��3 *1.Ukƹ�uC��|����8�y/��@��n ��j���_���]��)�����Q`���l6)/�q[@�2�AMU��i,��u�@|�_{#?~'���=�������;+�2^\�1bct!҃�8.�S[��؀i��*����ލ�v���D�RNۮ C��f��`L?{��/�������_��]a� (�����o�Y,���^�S5d�
��θ.��c��
���������<Ϲ�����t|�(�Y��X@x'��ٕ>�4���3��!}2�]�e��ߧ���}��o����_���ڶe�ڑqN�m
��4?��OY,<=9�k#m�	!�����;�|�q�M���/*�~`ڧL���~:ޏ��r��g    IDAT���x��	�}����T����_>�����9�����o�W�B�qxlH��뒗�`uc�h���'
�k\@�C	
��z���s�L2ж>z�lBǦ��1DI�W1�z�e0)�,��jr6lښB3�v�A�jE���_Ij?*x]NZ���a;g��w�Ok?����1����Ϝ��o��F4��]�igN��]V�y�^���]���_zc�G"PU{�<������Vk��?��˲*���
	�*�JQ	Ƙ׸n��������,�[�.����m+H$�Du�*���T�0�`�Y@w�5��l\���2r�:�D�����rd�՝�q��M�_|���a�ڶM��5�H���m0Nd�
Y�.h�0j_�~�/�x���]�ї���������_'��y���i��, �l^H�W^6~�v�@������[�U��{�ɓ'H/#���O��|����٬��2���&����#BE��%������O?;�Ó�G���/.iZ߳'��נI�f�+�(ڂ����\0�&'��j���10��|�Ij���P�%1��"'ONyzr�r���|NPX�j��dY*�I��  s��$ ����!JL���d�w�o�AVfUNV䈳h��+}��՟!���OQ��,[�B�e�QSg��1�N���^9?_�\%V��cFr��i��3�.3�J��,Q�.D2 uߵ��M@�v-�}fZ@,�f�,I�����B ���#2^������Cfh7�m?�i��1ﶰ���u߱�ױ�S"c�=�}q�����o�믿����׿�m�"BQ��Z�AИGW��ߏ�j��裏����Z��bv�W�q���B����a��M|�Dc u�<v�������U�o�u���N-[�y����:�su[_��&�aBiۖ���T�>{��������l�����|���ݞ���}�睛��Ƙd��4�8���W�s؍��k���|>�/�O�>e6��;w��?�c*�|��gt�S�9���*�M������/	�_ �Յ�m[...x�p���%u�����5�>�]�]������:��-QO[��.`]�Q��(�h�~��d������A��k3ʪ��o���]@>0.۟�4���k�P�=HR�e
�F�����d����([����&�Xr�&�&���_���<x���kpE�s9�1-U^2�U�U���1�_;bo/��9�+0���gR������Y��X��m[�������h�2}�=����̐)��i����o����>,^����#9U�c�Z��\�8<���o����w����m�K�~���\o�!�<�؈1?}�C���;8�����r���zï����j_W���<c�*�͆.���p�f��&���!G�`����7H�%K�A׶�8�������G�tL7XY�}9}���%ٗ8���� ��{x]Zvxn�����kw+la��4(��g��:i�h:Ď;�����1��Q��#6st"C�E��!�}�%���������L�b�f[��������%fk��4eq԰�g��ĎE��9��=!�(��?�I{�؝�v�� ����m[�>}:�F�g�`�1�F�:1�"�` ���H9[`l�f��X3�-�B��d�h�1l0����,^-j0J�5��ir��oY>=�,�4���~����}�EG�C����f�SBlh|�j�A�/����J&�e�/@
px�k��ڂ<? R�v�ɖ/u��7�^b\A�AME�w����,Ѯ�v-�2��A������f��g���~9ccN��9�+�l�D����%ưI��,�ܤ�0�1�brCk4Z�1ڦ���nr����bFפ GE��s�_���:�񂱞M��5�r���KU?@��<_|�>o�(6�>�l@�
��p��&Ȝ�7XSp�v�0�Ő�!(��D����φr�2+�v	�ѵ3j_�X��7��	��%F#y�g�>������'?ͪn�\�
(Lj�+�d�x�6o�s��|�����#��32W��!M$�>uGQO�"��
��hP��2a�˜�)MS��[�IZ���s8OC�Q�C�?C�>O�r�}%�
�:�d�b���IZ���d��to�|��>���|�,�z��<�ɭ#DM�(>��A�1�4M�E}��za�WEE��mOz}�z�K�fgq6I��2���uڶ�j����߼���|�?�����>{�����&s�����ͦ�+3��6t"񍯾z?~W�8la/�ce�|�FD�#�aA"���X�׉i�!�Eۚ��x핅R�EU�,3��JQ���Ij���O���اo����=�}�ݸñxј��#�m��دM#�ADݶ�4����G������u����E�/ұL����x�v�M ܾ6U�]}�0���W\_	=��k��9����Y�H}?SjS�퀚�ӅK��=� 2���y*�@���^�7��5j_��} 40��u��Q��,P���oB���P1� E�%��j�P٫22"��s|S��Yb�B�A'��5=���[Ӹ�=S5���c! A12�=���� b88ا����4vm��eܸ�*��������=��v�%ӂ��|�D�F%�U�K�K�["�.Y�Q��])Y8Ǭ,	]�z��,*Y��S�k�CQ� X�vM�58gp���}J ����M[?����b��n��;�?�=��&Fx������֍~��ۥ��eb�h�I��]��ד6\7�O������A�\S���\2 �ymZ�7�[_5�:����[���g5b1��ɡ9���Q�����7o�^{�����tE��˽�m�\_,�e6_/�U3�F��S#�]��߷}��oZ�����<�YQ�m��ں ����""��L�5��z��TkS�5�B�P�Fa6�spp���UUa����d��7��h�	;U��1[�U��&�]��U���tz��ƴ���s�D �l���=�Z�(��dw{���դI|��@z`���Ƌ�PI�{췟5�tL�8��ɳ�Ƨ��Ŝyf!�t�s�ӄ��D��	��:���*1�����CKQmϑ�#���Lc� &��o��Mz%VU�7c�����7߸����g�Y-ϒ�N,m���\�+'/��DC�$��{8�����oq��c��%��s�^�xM���.Ϙ-�S��$��yU�g�^�k�T���&}ڬ�ǿ��0�z}�����,�)���r���������#n�~��܁n�я��:��A�a�����7��Fb��	��J& ���4�b��%�EA����A4���;�dF��5��5upq�����`��uZ��"���Dv��a]�������$���+�͒��CL0Wҟ��cj��1q	p:�(�kDl���+��WOJ_o>�.��ʀ��D�����(} p��iX�ZxMר�m���AS;df�4n�2�޳W�Q�mӐK�yꮥ(
n�r��w���l��?��}���;˪�m��z��iV����xs1�F,D�R�ks��k�ߏ�⇻w����՘�T"�2WU��E����>-X��U��#"�,���V�#I�s�֭�a��a��i7����{fS�����Xh+��YFj�c�����/N߼<+�U�q�v�9Gx�04�쓼ܶC$qZ����4�t��)=���K���d:��}h%C��D��"}�Z�jV�����7g�<������әQ20eەί�>M�
27Ø��S�Q�d�lm�e	��{�Ǟ�S�ٜW_M�x�&U�&͕P-��!v�1��������'��G��O~��ݴ`,1
"I�Ӽ����v�dICi&�W^{���y��-�3r����ˋ�h&��U���;������<�.s4$�E�6��V$38��&,;H�-;���nY�qx��W����c*m�6V�Cn������َ��3~��_p~v�_o[f/��R����7��3�ԛ�f�D�C�;2��0b2��Q��!Y��� 6ptpȭ��̪��Wl6��I0b��XWR�,c"b<�j�!�b��eP��@Ҧ
C��T�#F�Ce$i+H,_���OÒ��jp�R�͘Aʰ6���6�S���ϧ��H���UZ�an�(����,i����ޭ��}�Âl��]H����9��1�M���s��}�3WV?��j]o]���~�)�g��wc�e�4*1�h�1��3k�ۨwZ��{��_�p�gf�����hL��Sj����^�MӠ>��ʲd�~��>�p6go��|���zk�x��#�:U����,�ެp�1�͈1�^��҃�ݔ\�BׯО��>㺆��k^�<wטy�V�<�����B�X�9�DljJ�2�y,�L}Ù�od�{ʪN#ik"\��DIiЈ����#��y��_9���#�ք����xd� 2�,2�5��%�cR��*���
4Kj[��� F|���[U!z�{�n�<���)~IYVW�EU�����w�Ƿ?�.�=���!?��O؄��ށ1U`�ʣw�1Ơ��YVp||��߾�뷎�Y^����?�A���31���f�7�88�KQkh�5{{{��-`0����O_	���`��㙼6-]<�����Yl����T`209yQ1�/8:�A����K)C1�9NZ[�1�2�~��F�f����g�c��g��,K�WԤ�cR��G�:^{�6��6�2G}@���K��ϓ$A��`�l$�8ź��<#/�5b�S�p�!���8���.
�ce��@�T�g�3�I�D�m�_�}�����W�����9�з̆������p.v37]wu�we?/Z�D�f.B?[I�碑е��,pրFnݼ��w���?;�</b�7���<+.���y>�WD1)�u�*6��uB��j>�z����~��G�_����S�}��_Z�;��9��yL���*2e�B�EA���w>��g%Gܺ�*��=���'�z�`j�P��{2��f��ގ���)=�|[�iD��1q���a��z� �E��)�ڦ@�x�=U%hD4�5�c�!�b^�bi�@���S{~�����Ę������׵!�������H�޸��������|�Wy�W�厧�����SX�3c뼘ͩf�"��e���2�8��r!�����im�y��_��[oP�
�6E�#H�>�׾hj_�GVV��TA<�ރ�ϷI4.�����⌣A>4�`]�S�%CUU,��KU1�3c�;��#J�6	��	�L� ���n6��c@���i6}���N�Pb��,m�+��;`V-�=m�4��u�Czw�L���8���F ���;䭷�Ҭ7|��4�ŇTt���8KQ��y�M���c���w��tmMY��Oy���V!.�J��,��&O����� ���#����QM�Z2l�0���P{�1p�����'�!�[�J[w�.��ldq��	�b	l��u`����|���5���W3�sS��i��U�Q|��/$�ug�hL�O5��O��{����(J�>9����N"q�}���Rڶ+˂�m��*xpV��hEPcqA� z;�����޽{'������~?�^�;==��i��<�L>#��W���1B�v���WF�$Z��#F�,fs||��|k3���X��\��|۷�I��C4U�%����*��]�]�qE,<a��c�^��{��o�
1�?ϓ�~(��7=Cd9���c��4�k��{���zI��&��F}[0��l^���&�9v?{�}���u� m�P�2I2v6��+\��Bf�TH$��9��R���$��,�c��;;�Ȅ�}�I�4-}FDȜŕe�X^\�֎�y2c���׷vm �P7�:��i���^�l6�(g�9#Ĉ5��o$��R��c:�^�8�,-�A���l:V�����-j��.x��"Y��Kתźl�oEl���4]ϔJ�K�~��1X1��IŚQ��|>6Mͦ	�Ͱ�@q��s7�����X���a�v��2��u����6
Yf�Ǽ��?���&�����%�M�k���Y-*���'|p�ۼr��1p��)���'����E��Nט�U��������v~���-��AŌڻ��h���m�R!��AcD#��Ohj75��B8�����j*n�IB�y�Wc���p���|
��ސ�麧����;D綝�ɑ�|�"�?;�Pb�Ȝasy�_���G�7o�8C[��O��������N��������w�<#s.�E�v!h�]�{�������㏟��~��ٟ��E#iܻw� ��?�?�P>��c�������R���q��I>:?��~���� �/��\������E���B��������ƍ�_{�;?ߗ��;NN��ƍ�z��}�}�������_�p��R88�{ĠbrUo��S���~t��òX�s�֫���u���s���G�D�z�O7�u��m�1��c?}nL�M������غ�z��������f��1P_��m��v|���lk����r�Z9]N���q"�5�ױ|��^t�v� ]��aHJ�^��	�5l\�!%�:�b�A7��Z�:v��k[T��4S=D�]���[Oȁ����{{{l6���3�,U��Q
8�]G�帬��H^�1���vKM���c-N����e�R E�M��,O��ITn�>X'���B$e� �Q�|ĊR��]�s�u	$���u��� z�w��	���kD$�����W:�ڵ��*�����t���mi�T�Q!
�W�=�x�=n��:o��O��qvvA�S�y�8�q�͛798z�7}Т|��O���gV���S�������MA�1�	���	D���TE�r2�0*D�
E�p/FM*��I)��Q�@��ԛ1�}��v��'#�&�gX�oȜܘ+ݛ�s�nM��� yW߷�^H
����7�րj�5�]S�b3�t�D�Ռ�����?���5~����������A_#OO��޸s��52�ϥ,�.��m�Vź��Z��e�H�T���_���|��;w�5 GG���%��������Ł�ϗ�$�I��O�	K�b�ң?�|_��������E��sa>`���ê�ͦ{s}e[�u�C��N���θ�+�r��23ޠ�>�O`��6\�����{pq�^�*��9�rpq�7n��­��m<�߿������߿��Yy ���9?7{'{�4M8�}*s���b������st�h���ߗ۷o�p~��G?x�Jl��[o������&ڼțu�:0b�*R�A:�����Z,�mZ.//q6�����.F888���z��7M}��Eu��l6ڶe�Zqzz:������*6�u]�V�Z����}��޴�j��}J��qΡ���r9�С�k Ä��y�f�T]Y�	��-��H9�HfӢ�uE�<��뚬�Fp0�G�3��E�,�g�u'�9��ֺ��m8n��� ��W`�"��U_}n�<�����()=��`�\ARu�b�@5�����:t��ia>�,g:�{M�]��D�#��o��2U�>@0`�M�L�R��:B�8���쒦IV2���N���l65y^��-�GĘ����C��7�u�|qH�>���:)��e�]�ڌ��QC@0.��L��օ@<1z��h�Z�XU%�YEa��B�ئgx�9��kW�hH�P�u-.�8#lV+�͚�zMD�7-�(P��@��*��Wdԝ��k��"v�h#1P��a}�V���xQ`T0y�KV-�z�Ū�����8���V
VB�$��ggm����5?����w���y��1mW��6MG״�9��l�ӧ?��<<�es�M�K�2����g3���8�.�H[7\�^p��w�N����999MծU�5>t=A�g5h)�=ڮ��"G������l�������Ӳ,�l6����u|���p��S��=��&۪]�����r�;��$]ښ�O��a=����2}l�Z�����m6���[�4��:}��|�T�b�mNOOx��o��W<�����=��������w�ʃ!{!���,�fM�̾��o�o�w'�?^���*Y�AbUZT���ܓN    IDATET�?tm�'���J�� Wu�ie�Xi��^D��5�w$�pb���ցD�x%8a>3�M��=Ʊ11ΈTs77̚�n�K�����;(Ķ��B̬�U~�l����n�cC�z1!�,����!�.j� ��<-��b\�}p�����y�ESA	������tvS�l�A��x�ez�7U�����N���6yfo��u�J��d�w�j���;�w�6y�m[h�7Z���E��f�eM����ʽPU��.+�B���W�;_����(��Vwſ���한��o�f�ݸ1��ixp||���������Kc��l6ݽ{�����NOO�\�5�+13Q�1b��ī��mT�n�,�x뭷p65Ä�&��׫x���(Hk�dbY�e��͆�O�r~~>�����:�Ŕ����S���޾)��g��1�u%�,��z��qS�X���)к�=F�>Ҵ-M���-Ӥ�k֯{q����n�~��b۔]�!b�	�5��8`zoH�5�0<����C_tS����`$1Y��a��5�-�RW��z�.��ζ�=�3�R��:V o{٦s�ި��*[L1DL��-$�kX�R�%M����#���p����� w۴ب��1U��3�;���,�łX���5��c��H:&�Ӵ.�)�j�6������pǤ�����g��M��)��W&y���i �@k��9���J�z�L-��J�U1�*M}��ܣk=?��g����|��R��s.�k���e�;ڮN�[��'�i�@����զtl"�b!�v��3��{�����3N>�9���}���;���Z��4�II�Ľ��>=y�_�Uj3���#.�c��̥-Cg��Q�˜�N�٩m��Bi�Ϝ�磌g�G'��4S��2�~��0�ͮ��kԍ7&U�Pׁ��u�<1�ܹ���G�����p��W8><B�ao��#O�HF��C����7����ˋ�VL�>е��T�C���\_���FI��Z�T$X�b�zb�eTD�Q%�kC1S�̚��D9��Β�J4)�*JĘ`����FUEĨ Q�	���V���ŒN�Һ�v��-&�L碪��r�ƺ`:�Y/�b�[G�FuAr��G�k�����R�h�4�t��D5��U�#&s���-vf6�"��"��\��3�f%q�\js�l�XjŬ�ܬ��;���K�ɨ8��1뎉�Hې�m^��q��q����v�7Y�B6��n6�ʲ�ks���b����7�g	٧]�uw��]��?�*��]��<W�$�6"#:rwӃ UUq���͹�\�&�ҋr��k����w���ZR����#...Fo��b��dL9�7Ֆ�����5ɼ2�N�=}�5�E�S6lH��_��_:��	�h�f#z�u�l6�Q�͚��s�����A#/��Tӹ�n��z�x ��(1M�:}��@H���\0k2��r��T[1�X�V���چ��X�X�8��t�2c,&�WR�)M�����B�5l�5���z�����'Ӱ��&{
��k��V��#Mo�������.��q����u8vb���4��L�"�u]ӵ5]S#�2G�;p=X	0wm_���
%*u����1X㈴ĘLq�
��i��8����₋�%��IkȺN�M�\"m[�&IF�u��S�r��[��g��k׬�K��a>K=�����Ԡ�>��Y�DB�@$������'_�����OL�5�\h�!lVAl9y���}�)Nj?������4�ҵB��@S�ԜG�rۉ�a�gg�|��߰٬x������O�tWto�����K=�-�؂:�I��ᗟӬ>�C]o�(�!y�7��#��LA�.H���yN����֚�|9�A�<�4ד)�{�� ���Sa���bI�<�ٌ�|��w���W_���^����6o��M����t1����l./8]y$*^��(���-2�yF"^���ω!��~�]����Uc�D��s�XH�D4@��QIii,�2�Ё�9�s�:^��X�V$��#U'`�%s���	䑪�m�UM�լJ��mG��/ۋ�.R��9��2�>7��Ġ��� �b{�U�:���;�մb��"�;�D�v�� �X���"�Y��Y�c]+F�j�1��m���a���F�"�=�EQ������i��sYQ,�z����ڍ*j�|]�<���_�9���e�֘�]ˋ%p�������������;�A_]ty��&hʠ��QTt��KF���IÓeI����X�ض�JFY�dY�GMI�W�%���G������<�5OUU�v5]׍�@�U�p|]yMY���8�U6oMi�i���Y���+����O�!�9��#��������M[P��<=;e�� �E��s`��:`�_"38v��A�b�^W$ld��WٶOz�4���ټ�xHYY�
�b�Tx;��I>���ϱB�z.�Ki��f�j���ҵ`���5l��?���c
=E,Q=b�X6�ߦ����H�3=XN��u�_�4�햳X�<�E�
_Hդ��(�Wk1
��X:�(�,+Fˌ�����O~�ӧOi}�f�b��LT�L,y,yQ�9*�xYg&Q]Had��������euq�/?��Y��3�g�,�5�I�~���)0��)_��>?��g|��_�o�;X̚�fɬܣ��j��_�C��/~�j�%_��m�@�`G�/"��Y��1F�&�8C�����˧���D����%��4W�A�8��2�|�!�D�"��߰<�P��9O�dY��U��!ec��~���y�� ՙv����{�n��c�_�6c�7����fX���dY/������o��ݻwy��w���;ܺu��2+J=z�f����������U���3�\�XV��lV�Xra��QCX��^���������Z??F�у���A�#��p�$1���hLMf2p��b���Q�_�W��!QP�H��QM^���9Y��ۜu�f�L��b����d�y�'K&�I.b2�JW���^ٴB0�"�)�N~��)�C�tmMYU�Z����QU3k��]�*s�͜u��1#��ط��?~}�f0ԛU�%d�r�]�|��c�Y��ږ�Q��W�f�Uf�jU����5��6���lfT�s�޽���/�l�ݻ�߻w�u Gu�LUz+f%BkĄ�D��$]�GP�\^^0��{V.5Zo�^�=UU�h�.�T�1z�>=���?�����o�4h�|�Z�z�M��=O�4�cl��vZmE��=�wB�� �nzy:AL��>��%Q���j�����jE�n�,/Y�V	��X|M`�<�7�+���2��1���ܚ
�5J�"5�u�=����!ڱ'��@4[K"�B�'�hVL��B������:�e;QJ��뼠�r2�h75�J�:b�p`ˎ�L���mQ0���勉�7��q���l��2�U�@LbOڶ��Ռ�#�����T�ٵ=�*F;Mc�j��ɖ4y��r��|�.�s��N��g?��䄳�?9�r�ĺ2u����9\��l�TC�^D�C_v�7ہ*����C>���'>C��e)����zY#d�u�1zbH�e-g��V,O��~Uc�ʉ�MK׮Yy��?��_��9G�ѐz��%EL�O�4�}
�<�F��<!��q���"��!u�5	XxLH�%F�@�,�-�� �ΧjQ��Q�1���t����3�������삾�rw��s�f��;�i1�n5���0v�߰�4M3j\��eYr���ַ�Ň~ȝ;wx������S�5'''<y��#'''<}�$IDbd^Udα��鹱�!����S��l"\��Ҵ�����s�ME����h�@HO�Q����'�*4>��:��#t�x�Z�HD4�&U���b�E�o���65��3��_�w�@V�bFUT	M��3��g�+	VEQfe���-���(������6_����w��	IA��-�K�f���]��B�AIsL�<Yn������9(ɒ�,
��84up�\��ǒi}�P_�Y���(1!�����ˈF���,��6�1�%��T�o����;u~����'����2zF��1ƫ�
	�mu�� �Ba-��E�et]Cy���z��Wcx���O?��Ǐ���P�8�A�T��\1J��tW�)?l�Tp;�wx}�����@�n:z؎�x�뇱��M�1�"�	1|�5��6��כ���r�Rt�b~I�;�M������a���6���k$�)�#^=�E�<g���J�M���\����V��CϘ��9g6�(���,Y.�����L[��:�+d�$1}V�zk�:�˔��6�Ib�D��A�4(W��q��A%bI��vQSM�Rg�������ᕛ7�_�Y��ҮVtю۩�	�����٘��,x��|����x�����!�͆��'�כ��i+��a��rA��1h20F�$]c:{d ���EAS.�fţ/�8y�����e�6�;3���C숱E	l��B!s�e��
�Ո˓UKpdF(r��j��X9g1��3L��&}3@DL�'�TS��JJ�9k�3A�@7�ov� A����JJGG�(iaF�,�e��Yb@b?���oۧx��9�g
�^~��n����fC����9oÜ;�����zF^7���a�If�u�W^�|�=n߾͍7!����>}������
>65��2��b��mq.�陼���e�q�&����1a�*��Ҳ}\z���ɶ
��t�-��ߢ��]��X	��q�$�g]�X�㚀!1���^�Q0�.��M�vE�>I>���l���׈��9�y�&��1cG�$ˠ���R�r���ɈJ u��yF�2��T�%�,f9�2cP�X�O��h�(+9�
K�}_f���l��|�N�1l��HJ�u�
E1��m!���9B�9���w�m �#��*���f�[%Rh�)�[���Kg�����7��w�����Y��k���άx�������N����������0ܼy8���g�<�mkNN������/��p���[am�6W�����s.//��`)B�� �)?ܘ�"��=�vR�C�7����ԎcwB�J��w������x�i/d_��,i�+��~ۺ��/;�=��{�{~�GR3���<�Ry�[6��V�`�6�O5�@:z4
y^��w�|V���M��-Ѥ~��& 7'C0Q�%7n�^�7nQO�<%����21��~���p�$M�V��h�5�Ѻ������,�Y�\'����C:�,
n�����Y-988�ެ҄�@�Oo�Q�$�#�{�=�~���{ұ����$�1E(-i1r����ʶ�r�?��'Sˏ���muM�u�[%�k�h�v�#OA`�2fW�$��X�HP:�P:a��G�u��k\!�'Ѡ�2wX�<��AN�Z�]�cj1�ơ:y+�u��H,t��(���Pa�$pb��A;\JBh�cRP#�}�qH3�y_̐�}^���~�+�kwG�7���u=ʑRox3�q�5e����7��{wg~懁�\����|�[��7��1��'D���3�e7�u?7m�]�B�D��XI�<�Ec�n��J���Df�\N�k����{'�="�:��ύq���e����Σ$#�:4B<6sxBj� 6��GZߑ�> �B*�I�#Ĉȝ�� �@��f�X!w�Xd�e�0E�Yr�a3�3��f1��t\� A!*]���:�}�5����.�t͊ns��| Đ�m�~���@^D���C�v[>��������:L�UU5� ���p�Х�S�3�/f][w��NC좏A�uU+մ���<��o�7��o���%��+������8���w��l��d��[�$˲dnC@Fd���h�Q!�4��Z@��4�Y�H��;�l+��lQdS$��*��>��{�W�����[,6�d�[\��{��s����������:3Ea����+��V��pe��$�*���6M�Ǫ�B)��#rt�<R�nx��>[�=���bI�?����G���`�e2�\.Y,}szk-��m���1m۲X��*�d��n���tQ�"���X�'ɓ���ٳ���/=�OS[j����%�"*>�inO�7��8��V+�QFf�$����c�Y s������{�?�'龒/��M��E�/]�D�:}�8�X.�ƚ⌣����^~�+7o��(�{�n'G4�5���ڹҝ�q��2v�PQ���y����-�w�,�K����R�J�㒋/b� >��3��T��v��Z�b4�=s��M^}�U�I�T5�Uloo�2��H�Ef�Hy*�1����-ٙVYgm :��m�7hi��[��� �!A"J֕�:E_T\��ʁ	ˣ9uh��꺽tr>�1�>t�!aRf���P!�+|�$��&֩O�Q�' ��������1:�I<Zi�*pc/v�`��v4�%t�U��6Fw�����E�c�>��
�g�&�;#$�EQ�sz�|��g{q|�kG���u��7"���+wS`$���Ʉ���hc*r��f�6@r ��>�9:����@T'	�x4�{߯��<���(ǔ�s�}��yR�Խ)�&b �،Q��I�Q��y/$"X�is
(��z�����fٴ�I�ת����K�M��p&�&t�=�x���m�#�Yg�T��x���!�5e�h��LG kM�mn�t�kޣ�f6_���Uv>�;�+�R��&9�J@ɺ�(ݣDq�����z��=)8(�(�Qh�O
o�|�4N���m��ku�g%)�b�7��v�g����y8���6�`�\n�j��R�a�VƳ
�� �ˣvw/���G�������oE��W��cV͌�?�1<�i�Q���NgGL�SƓ�
SJq��5���o1����8>>E)�1ާ���½C�^z�� O��4��S݀�<��M<M
k�|/����~�w�|MӰ���Ç��U��H�>Csr�À
��D���dZ��-"��c��e��e�x�����I(���ւ�&�Ef*xT�γQ&j�)>�B�&�:}�_�w��g`�g����*?EP�����Ũ1Z�)ѡ�Q84���*��U��u��	%,������� �#C�u=�t��&E>��[(�͕K/s��_���i�@�\���V�d-[eƃ�Q��'(}�>к���Ӵ�n	��V���r�EE^��$��'�a�jE�F��<�,6h2Q��튑��Tx�Ȳ��Qň���k�����OJ����]v������������#��=Gh�dh�O�=��l��K/p��7(��x�-��'ӆ��.��㼦�9:�,��� �
r��!U�nF�d��	8:�E ����ۼ~��ϗ^�1�VGp`u�!J�b�fg?���},�cE�� 0�.����%�	�Z,G�n
13��$lN���.�$	��1�����R"T�l^;�B��0�D����9�=�E)��!�t��Xaӱ]G<��iC�,�Z�3KE�6�M�~�a&�5m� �-�uEU�(��_���{ h�(�	�̡E�#}(pz�b:ً �$X����h�K��B8�+\]Q-��nUL9��<\���1h(��rdg]&J�>Z��fvtS��f��"���,�K�0:��y$�Fk���A��W��9�w=H.�H)Q�vx�����������c�AE
��cg��\W`��|ۯ��1d���sWW� �#m��s�(�ƪX���=H��#t�_�����t�������ޭy�!�u0�w bj��߭�Xkh3EU�m�〻@�n���
���g^��V>�˗������,����QZK�����/�M3k��f.�,��[���X���~[^{�TGs�:Q&[��G =�/^00R����]�ܹ�������l�����[oq��-����s����}�:y\GG3._�L��ܹs��x�o��o������1��ǜ��Fo�5�D�>�mvAaRl?������3Q��%�q�<�x��ώ�������A��/y�q�$ �g͆)���Ǒ�i��p�N$����˼��>���~��l��tL����nT�%�h¨�H��]���Q$ت!�    IDAT���ZK�t�g,΋&�s�
�����cn����I�$(��	�������C������w���s�Έw�����M�v\'7�g�$�j�(��4�(��mFcW�&�#U�f�e?�lΡ��t��j"1=�N/�E})���9�Ʉ�,��f(5�����⠦*ߴ�TŞ@�s�b,�E�&�u5M�hh�S�ȳ2�.���G�{��K��c��9�u����1%�^kF�6��!���v^��6� h��^�0�D�[���B����c!C�{T3�H}��#s�og���^i��A�1�����k͙�cHAm�ޟ��M_�Sy<�;�:Q�E1>�Q޸����sM���.�����m	N�:C�eUD��kc���7�o<J"�w�d�e$�v��܋�8�*ˊpp|�����w
�G �������?�C�]��޼Y��� �k��R��cVr�pV�>��5�����.�"G#4Պ�Ǐ����������Xr,QH#��R���n:����)z�"rC�B�*|�=o$i�����t�J���l
��0:8l�A��c�{��QA�<��8h�Fbi��l������,[�xz�*����rU�ZF�͛7��sz:��dƅ��Oڻ���uǁ�vc�w��^p.��<�êm�yG���?�����!��LS9J�H���ˎ�prr����v&ܼy������i�k[�	�CL���E�<����� ���#tabׇS8��Q�t\��6�{?c�o��yLrf<�����>�eY��|��QJWN�v`����D��<��g�1�Z6t��-�SB�ڵ����"h����ƍ�@�bQ�B��Oiac����u�u������i\gl�G0�5=�xPg�ADȳ���E�����Qx\��u:��Е�F]>m#�/�QVG�<4�9B8+~�;�f�A*���,������"Q= �MA�������ߪ;��<�FY��:��˝t��$f�b1�CY���F���mQ�>q͆�2+#�,�."�u�w��Y�ʺk�#73�U2B�m�Z�"�����o���j9�EaQ"���m���ҕ�!�6C@+����޵�Z���K�$�E�G�j�/!:h�1�`D�&`\��YU.\����;w�0��1�0�y��1"���1���K$�:����������'�'�y�7����aLy�/ے��CO�i���Mj=_�[�B���Ң:�H�{�����s�>R
$�u�Dzr������.z�7�{�5i}���{�|>����u�L��P!`MI�QAp��l	jF�j�Ν:�<~����ׂ��3.�paY���`�ym��\���s^ʳ�~wi-�c�����e���)M2.^��d2��e��:FZ��!�����f\F3���� &C�"+�vDլhR�����I�����>[�-�Zk泓/|�Cg9��ZF��ɄK�.���)B���w������D~ga��$�`�eU5� l��q��M�]��x<a:��X,9::���������+ ��M�^���3PQ4f��<���Ǒ�qڲ�k�ީ )5��1�'���(���҈�B'���X|P��<%����FcTWr���+�Gi�o�t����Q�%η��b�Z|PH��wxӤ1K �.E��&�4!X�b�������L��@b��&�,�z]�s:�E�.j9�?e�"�v8w�E����z݂5����G먣���UyL�g�}�I��EiqU̈�m��AME����V��Ѹ�W�9�ۣ�3�#�[��w^x�;��*S��sJ렻�k:r+
��'���{�6Mӟ��Ǐ{��h4:3�����t:�,�� \��q��3@+=\=PROO�~�J�{I�A�.���K��	`(�YeY��ks�9�=˪�"�@�QJ�R%�D>�ha]������'���&�,��$��v�������>�d�A9������~x�ӓ9[�����Q�)G6��E�ꆦ�c�$z���wTZ�z�ꊐ�wݤ"=Y��l(O�"���2��ֺײL �L�4��	=�{>�s������^�ҥKL&��S7B�:ڦ�Y�>�>�t���kb�m{{mjZ�ԡAw"��r��k���5�yub~�l���X�go�y����km ���ŋdY���Q/���Q�����Y�ك���O ̘��vQ�ƹ��Zr��n�x������3�{~kh[χw�X�8::���CNO�q.tѯQ&��:��d�h�Y�#%��E�b�61���T�[�4�o%��p(/��^TҴ�V�d�H�Ġ�{A;���(c��|���V�C��DmE�AD)�h|z)�D;�Ĉ��:u唏Jv�p��w������N��|'����	^�(�g��A�V���V.x	�uo&j�k��@�j� �R38F%�{q1L�<*"U!T�~QJ�6fuナ\� ��AwaU �e��Z�R!�(o��D�;g���5�5���7�m�Ci�^���~,"�d��cT�#c�_TҾ$J��.���D����+�>��ݰ���p73jn0�AS*��.�b�\�΍�e�|���I��h�?$�D�;���ӓ������dIѮaĦ���q�@�{�8�É,�8�ӳD`��ϥ�0�Coq��U^c�!S�p��'-|�&���`C��� D�D��mt6Fk������H]��{;���(�mmAS�hcQ6G)��9Y�DӇ��w'��gr����y�g�)�ϸ�O�cl3
� +��5�c��tM]S�Z��>����6#�
�wH먛��ZRU9M�p��iA	YQ��w��tBF���
��h���D�6��	"���f�yk8&���:cl����(Pb�nR�T��g�\��ߟ�'���kU��7�=/��uv���F#�˚{��������x����rA�BuC��y�Q摧�"�Q�b������x\�}������4.���*���.�j)�̓+�U�#�#"!��˃3�6�B������Ҳ����T��SA\�ֵGG{˽�����RY�}���De�5~���Yf-#�m0bt�G^S*t���8��ʊ�hU(��X�j��)�&JFi�%'�$=�L����z�u�M�h%:+�P�X<+�m;�����E0
e�Z�VDƙ!H U)%�U�P"�(gă2h���H�2�J��A�ZKP��֡PblP%�5�eZk/F0FBQ0� ^,J�,ӡm�>��Z���Ѫ��ӣ��2V�8����Ց����Z[?�,܍�dr�v��}�Mu���Fo�컂:2YvA!c"�[3�6�\p�ek:��Gwh��o�@�4<~���>ƌ�q���0Ĩ�V�>���9�ٌ�ju�T~a8mxF�睴��lP���P�~pm����I��a��a$q��F16�_�K�mʒ������OZ��l�D�(��f$@G~L/S�����M�w���{����d��$[����f��ݝ��&v�(�y^c2�9��}�ш�h�<� ��{�6���Kkr�9�{Q1kL�oK�hkk��ׯ������#<xR��0x��������-�|�2�Q��|�ֆ�V������=:�{��p^��+{>��3M���%��-t�R���u�z�g���I��'������m&*���>^�o��;o�����!��
�'�:[W��6��&F)3Ma.\�!/3&[1[���y�_�4.��yh�Z{�B+�.�������v����+���b�ֈ4���MF;�V�΍��b]v�4�,���R�UVm��.��x5*���3����o���_��Q����O�(�~�w~'�����z���۷��۷�J��}�������t��6f��R�c�ƹ�Nm�k��f`�UJ����{�L0�k� w�X�TN�h�>�,�*����*��\#�l�:d@�dNkk�C�Pʪ�����D9���s6h��Z���8��1GΙ\i��֫;T�+��*��Q=��Tv$Y�a0fi�ʴ
�m_���AV%e����t��r)�nݺ%���8��Ng�ڪ9Ɋq�> �Qd���Ն�ka�X�e{{{����������wI�(�F��szz���J)f�Y�oW��x|��ؒ,�đ�`f(�.�O�g"��?M6��w�Xd��3�9�ߔ~;����6
9λ?�`/�ֺKu@���Q�1ژNGS�N���}�o��_W4�Q�Sc3��N2�����۟Rv�q6/�F�	�������g?�R��|Ч�O�*;����"`C�+��˶��ӊ<˹|�ba�Px����b�xd���ĭ�H�{)6gw��l;�T���k��
5��Q��싷D�I4X��"�T�2�s��Ms��x|����ŋH�O���$SJ��|��z<���ϕ+W����㣏�����hm�K���!f�(W�5ň�t�h4�����x�R��|�jYc����\�x���s�}ur|��T�Tm+�r~$J���EU��AB0^���ki���Z{�6M�hT��f��*��F���fbmc��Bp&��[���=���mk�x��znL���҅������ (
;�sY6��۳���ܵE]x_Ε�lQd�z��������ʭ�n�ɤ�>�����7.2�im������ڋo��}���X?��P���M��,�q�X\�U0�h�[��º���(-
_�F�bE1c\��s����H���Y�H�@��X�\ �i��~fA+������ked$^��z�DNuΞ�m�>
5��⼘V�4�B��ʚQ�C}\Uvvv�yؒ�upppr��α������p#��TL����0S� ̛Z�(T���;��{���_����QJz�w����ۿ�ۏ�.��o�b\������-�7�#����"3�l�o�V�u��+˲�%�#�u��UJQ�%�ժo�^�6=����CUU�C��]�Uz^�^� ��� �
+��<Ŵ�a��@Z�=��E��(h۶��=L��57'�=��x�5Z"6U��^��%���15J�v��Uk�8����F����f�~Y�(�δ�Icዖ�I��kK��g|��f�=e2��)�4� ����	tc� 7e���Q\�ckk�+W�2�-K	䅉�]%�/E�Z�p���^<�|��ޅ�4����qɲ]��~�yE����bу�ƹ56�<�_���ñ�RcQX:�#�����m-��˿��_������}�փ��gJ�G��:g��*>��ӣWؾfI�u�f�b{w��w�f�4��X�������ϊsǺ�?Q/"�0F$�#1p�6���~Y��}=+���:�_����ܴ�j�Y]�MK|��y9͛OK����,��y�h ��^�\�l�e9�aݖ1uu�	����Ɍ%���;�$x�ݽmnܼ����'�����&��"0�n�H�R�՝͉�c,Yf���t�r��������a6�ك�G,���nX>>���cw�?�^�tq�T�#4{2s�}\�֞�.���i''ƴ�͛�	ʨ�6�������o-���\X�.��_�z����)��śo�)Wo�R@�}��p��������խ[�$��?�?���۷��q[����i�[�n��&��81��G�p�_v��|{�j�]��6׏.�ӫ�h�ԓ�AƩ���q+���������cK/n���T`��v�%;ń-�VK���YQ�e�L���Q�y���*7�(9����ж���8�Zoy�m�*�B�h�5tЂ<��h�WZ�v��o��.m�z�o�����t>����Z!�F{��2�����R&��y{4�O��T���O�a���_[��{�;�V�daU�em��j�7�~���P�h��L_nr!��4;/�;�NY��ʟ���j�t�Y���9���
'''����^k:�TB~�bك'�؆*	;'�2�ȟeK��	Зe�d2������O��[C~Q�����$o�sBw�ӭ>*����(3�>���u��h�B���Og��Ιυ�����|o�"�/_�j>D��Gk���}Ї������/�&t��|}���-���:��p(C��2�d���|������obm�\����w?���lxZ����Z>�w����������E��@v�.����1&>G����Z��OKe�Ά��������$���s�k�d����!t����p!"�����8�
�>�E�;ֻ��x�y�w89��M�@u��Hj�f��s��e����L&�y.Jf���?�c�֎�jI�liZ��DJ��X���/�)F�����rn"A���eL���M�����?�c� Z�Y/9�o�������7���|����}�7��称$���R�����۷o���}��Pr��n�|�p��5�����0|�ߔݺõ�b�r�ܿ~]F���|�W���C��pl ���t���N�>��ӝS٫���Ω:9��s6|��U���?s������y��ξw橺}��o����<�Gʚ�b�]���՞Blh%7Zc�A�`}�&`��k�h��k�w�F<�����-`��rN$h��$�L5}R�i8qE��QL^�P�15�NQ������������2C��tLÔ���kj���gV�ՙj�/Þ��?��he�dfY�Ot_��=�6�
8[nm�F�hm�6�茠3�����ϫ���믿��䐏��ؠ� ig�OS�𐃇�88>b{k�";�\�|��/���Ǐ1&���*�;ϔRԝZ{��t�H|��<�w^Tf�K�u�M�(�J��/�"��k�dgg�����?�0�y/8�e@�v�w�i��"g{� �/���׏�墦i<u�X,*���"����Odϊ�mF�����?�g�<ǻ���p�ĭ�4B�]���o�7�����������|7�4�`�Z�4v��4k���QOK�k�d2�{��f38==U���qۺFIl���E����p:���	�R֒�F������iZ�����~0|_YgO�ގ��O�?z��I����g�������+���%s��<�ƨ�J�C����R)2�Q�Z�c��nMQ�aUk��eC;�K?�;ϔR]A�Y��M0��)B7�L��<�{^�d2��ݻ�W6L��xs�J�F���1G_��tނ�,��������%����Z�96���4�*��E�X������|�/���������گr��>����U�B�3���̎�m�v���1<~t�������`w�W.�@fe]l�w�OM)n�Ϳ���i`o�vFg��YG���d{o��f����~�G���9M�8�ɰy�V�K�>��ݻ��ҋ\�V���u7��d�b��,+O𚂍9dy�Y ~��=o�w����ڜS�c�,J۴0P*n{8o?������4�V+NNN��&���cҧ]�γ���
���CB�y���h΂�$ӚR�%�{i۶�C���'�h1����g(,J.�c�Wa�X�Z��d��3<R{q6�^�ܮ����m���৛��ʾ4{�]�������r��ҏ�׳�LByn��+q���J�]2�c�$�`:O{_Q� k�6�Ki�a�5�!P��_.����V+����,y��^���i�i�3�жѻLಪ�/�����yD��'"}S��z�I�y-ݯ3i�n<E'%�)�����C2��6.\�7�7�������_��`�b9c����g��aC�����֭��؞��۾��9��Q�m싊���o���y�/����`��˛�g�=sJAQ�i}�,snܸ��70�PN�������o�X,��#�#vDц�4e��ʐ����#>��C2{�����or��/]�i�?�׊�d�	J������m��l)�5���ߟi���cꪔ։��e���\9
|^��M��2<uS�C��4��?+�w68��{�ɘ��^P�X�����Ƭ���Y��3�ǣޑv��Ѩ�(��Չ��RH7g��hC�EY���2�2U(�[�!s^�9���+�[b�&n��xG�2[��X	�f�F��|�t�Z)b;�4 7���;�"d�҃�"�	��7�<ͳ�\7ӥ�{m��)�ato�In�tC,�3&�oP)�w	FiA�.    IDATӾ7�߰(%�y7���h;oR�=+���Y��t�S4�y�3��m�c)�O)E7���Y���7n����_g:���ጻ����!YfP��9(-X�	ƠuL�<z��*ߡ^�ܿ�|���'�FP%����;�?��7ql����.��9[�z#}��4M�`y��5~����|�"Vû?>������?��>~�̒)�hd�@��Sa�Ay�.�?�����-9x|��l�h4�,&�W(,Zٙ����7�=o�����p���,����9t��Na����f��y�O��l:��U��c�ٌ�ry&��|<��[k��f}�.�S�EQ�Y;����4���c�t�I<�bKw��'`��G~�24MMTԳ4�w>2A�w����n��~�\�W�sjO��۷o�����!�V��^�6<ԙ�����iM�7Z��(5&�Ch�p�I`( �1*6D�]oǓ���dO{�Ҥ��KO�WaO�o��H�Q�}��[)�Wo��䱹X�m�^O0���,��Eq���ާ�__��霡�7k�N��p.6d�&��O��^Rᣏ>���j5�YΩ��Ѹ@���V�k5�讗��Ǉ8_��c��X�>�YE���t�U��F����ؤ(el�A*�\t�3 �<�T��F��OkM[�k����h�[o�xp�.o��gܿ�6����N,�<뜥��tJ2Z�@k�.62OQ�?�˟��g<f�#��P�<'�3$(��i��r�i87�\W���6���������O�<?3G� @KmS=1ߧ�|E`������t�S6g<#"=��yl�����ޡX� �@p�.�F��J89>\GJ�fT���m��bբ�� �
�VC%
Oӈ4M�
�[�L�Q���vF�90����)����,ٹ�Q�])k3/.��Pg�}O���J�Q!`�����d�ė�b�C/FDX���Drvayz���8�D�6��":	�=�Xy����XP�0�����0�;�,�g�����E)�{iC�/Ҟ�>P6��I�NW�ŧZ&"]�óܸ4�b���µt�)�lmm���͏~�#�̀��oO�u�B�Z�� �Y����s���|q�X�W��bww�</�>�is*g�>��,�"{���oq�ٟz�r7>7�8&�	����~������7?�G�<E�S������kY�jl&��S�(�w���ȩ�#���ׯ_�������cr���?�B���3�u���
�}
�S)c��E�R}TjHU9�c�4J�$@5�N�N��-e�Ζ$��|>�[�����9�a�#�L�,���<U�9���L��s��i�_k���.�l����YUUvMJk����s����s����S���i����Yn�	M���Z��nf�}��>z�b���g��}������~5b�߹2��������B����4���]�[�Xm0��j�kO#^<"�F���-1�:*yV���U�j)�:�������kc����<�ŝ��j�a� .�u ��􈭭-��'��R�5Vk��8�Hal���m��2�=H�w����
)LqH^e�Mn���� ��7����0�>�i=�d!�I}}4J�j�r ��/h��>��� �8�ٚ쓛-�Q��&4\���G�,���;�2C9�?~Ŀ{��</��?<,
l�i١�u���/��ͪ�����7�������]>:XB�^�ԒǇf^�ƉB5�,���	�v�-7a��<^=�n�r˪
 ��Ni���g_�O�JYT�G.��R�j>CG�ۓ4C��j��j��
5���|�Ο>)�n����F��j9��Rж5Yn�ti�w����?�x睿���nG<<<��m#���B>�3���sC�t4M���1���$m<��=3(�S�Q��ի�2�@�C���D�z�jǣW-A��8��*�0�,���S�4ԋ9�լ�m
<��&�B�0
�P�סu���in��]�������傼(#y�	�B�`	m�$p��un\����.{��\��C�@�\��T�GǏx��!����v��Op��K�0s-��2�C�U%˓%EQ����o�̅+���,�(Ǹ���vI�.��ӓ����]��>��	�r�xOfGhM�'�ھ�Py=�k���<!�E��W>�Q����1��h�s�����a:����@�E��<��IAr(�����@C���-J �Q�f�aœ�����Jk��y��"u���N���Zw����P����xoG�z����Bi�l�������WK7�������O���~��\���o���=�2f>.���j��^cj����5֢۞ �4C~�Zb��^P	��k3D�D�C���Z�x�}�6ӌ�s���\��e�G6�|J�*�,�X,,f�u]������"ҡ� n� V���(Sqq={��@Қ�xn���m3f�%J��Ձ�N���E^���SLE����Ÿkf�Tt(��歚Nݿm[=���½{�x��8<<�Q�=��hU�V�cMp:>'*�d*�x|h#�V!v�t��QT֩<?;�ƒ�%Fg�ҢM��nɣ�����)A��Ϣ��o3M)�	����߽�|�[����V@��ҁb�T��}�"	���"Q�B�M4����{���(���X,���u��^`o\P��`��9_�3�/m�B\�t�Wn\���q+�ݿÝ��`��j(EfKP��n"�����y���y������&�g�2�h%T�mUst��;����ŝ�����4%(KnZ%,]|V��x'x߲XԼ�����_����Wٿ��YD7�x�i��+����f4.�t���O���(�5�J��by��<�j��ß��ݼW�"��66i=ß�s����q�7�g���3���y�X�VH:x%X��"�y�T"�{�ӗY�ʾT;�����w�w�R��j]XV�f�ng6�&
�ɛ8I�c����'GqR�s�s)-���#�=@���
��k#�>����,A{�Ɉ\�OJ����ސ��Ep�6�DHN���x�ŋ�����?11}��������*bH�D%@�z.�����M��"�i�g4)Ȋ��������A+E�6<>����9	
c�و<O|��H=��aZ�1���,�Պ���>"�:�y�5
�"�4�AO^(l�vEۮ�"A;R"@z�;x�"�@��1�"(�r���+��w9\T,jG��,��UZE�a���go�c�a�~W<�bXձ��6�ۮH�K�� �G�b�QxeQ0Oy�k/�5E� �N����� l��2���ɚ�y����y�+��/�2�ܼ��*��>b1?��g���2d��ʫ����_�����^���S�?z�S-�q���-m�	W.]�՗�ί�����.��۱���)Ah]C>�c4Q�w���^fz�
[��x�wx��~��f��[�LV /�g/�t��|�;|���foo����и��ű� �5�0��^�0#���������;�NN��PZ�q�i7u�L�9�)���?�o��͹<�p�t�a�es�ߔ��<��-��=�:쬳XA���������n�h��X�쩒���X���$��|��Ai��u���kk�1z�m�A�A	��Q8g�u�IWu�G)Aa	�j��;#��^��<'���R�^a�Le>˞
��0���,)ҧ�ꏡ(
F���詀��MЗ������C�}q�TmC�^^��#��.b
��e����%`��Y�,�Ե4��j���Y��������������hM�+DJ�(�#]a��6Ɠ���5M��iWx�PZ�Fx�vh1���6*�"|�Y�"���`���~�%����:�V��h�Q�z[(�� �Ƣ�b�d4B�15�X�Ed5>�h��]L�J�Պڭ�m�����h[b�a�j����7��˯p���fww7F�f�UL�F :-��ŗ`"IX{0?)�6�[��ï�������������d>;��Š�k�< ��1Fs�����7��.�v�l9c��Ĭ:F���-uAqq����_�W�W���+��&�^@p��r/�����/��7v(&Q�6*�����T�C���8/�G�ܸ����	W/\fog	-u�6��и�v9��
�������gS��0.�@��f'BL�~��Ր��C����E�Σ�9����S@�y������y�o�3�u��:�"H�v�!�J@9	�&�p��͚�~����?����o�=��1Yݢ�Jk�k�2c�dJ�1F4�#)��#h!�yDp.����ćF��Ak,��`i��0x�o�x � 7�~'��>�ڞ�4]c	Lӿ�ņ�J��$�Vp���{�r���Çgdl6���P�ŚD����F�I�9��9Z�Bق����Q�y���Kr���LIKp��b^��(���2��5���D�5dV����P�U{���J)���L�#7��ޔk�.q��.���|M�V�m�-YG��#�炀����F��4��1P�kF�l��/q�i�Nv8||����U�����,Fi�����(�mc�⪉�������zE�j2cMs�<��CPh�c���=Ⅻ�^����J��y��&���Q)eh�Z#�}����X�<�(A�`�G�B���/���OQ�(�c����X���~�ݷ��|4���m(Fc�|L�!
��,˹v�*�x������%���K<ZTg���%�k9��|7���)�\�V���3޽JZ�|t�YՐ#P9�5��������^~�reP
��������G�G�mC����/39�Ɉݝ�}��Qd}��J��ɊŲ��ʀB�|����v�{Ӝ�Y��>;�^�y�\<�T?�ZO��͵j��u����ӂɩ\��UW葧�� J�	��ҥ����9���SA�t��
?E�Z+'(U�km�3�kl0J�lv&2`�A$j�:�����K�$Yz����9����wuW?���ְ���%��� �=;o	A� -�!�` pe�2�YX^p�	�m@/J�!��GwOO�����Uu�73#��yq�䍛uoU7��d��
�73#22"�9�������-�@���:�Օ�1�Cx���Y��QL�~Ƹ~��#-k1N��_�����Q�ũ��l�<����9�#��:��?�������C'����#b�H�KPK9�������X.��)�E�`)�
c�we��'%��s��rs��Qb����I��.m�0�l0T�0��h4�Kk˽�q�˗np��y��g����7�d���_]�J>����EL����I�=J}qcs��|�p�ڳ)�8D��'�]���gOJY���ރF�g�J�i�PVfU�j�X�P�:b0����U�=��te��J��bZ����3 �g�N_�S�&0m��\�h4��2�3JYV�;����7���J�RVc�rD�=��PE1��¸������3����u~�������rI�l�}�}>���N7א���a
�_�t�+W�����-`�\����K�ˇL���/�����+��ʷ��[��)�o}��������98�vc���/"EQ�������y���v��8��mv/^e����]���"�)}�qWb���K�
ﮏ�}w���y��������z�����ѩ�ߕ�;zdH6W�"bQUU4�Z5z4n(ԟ����s�ν؛��Z/��}a��3co�m�s�)�(��9��t��J���w6 5mk��E�D�K���H�1�`�0,+$*N�%��@�Ā3��Y�!>d��Ͼ���\w�㶼�<��C�GGG�t�<�f0�߶���&�Riׁ��`��m���FM�%�sn�s�����J�}�l�Mݲ���ݻ{�
;��xV�.]۬�	+Ч��iq ���KBlq�d<�Q8<�5���8�M�֭�%.^��d���&��$�C�E�jf��>�I��"R�c&�{�
�VL6�lo]F�"QY��n�,����QU
SR�I���RU����!��h �jD
���\��<>�2������������Z�����M|���>{g��I"Q��;��u��-��Q��5X�OKA�C%�
'a����}��6��!"W�6D"1%�p��3�ʯ�:������K������O�џ�	��G?���vl2�.js��5�?�W�^��SOq��5F�1bK6����"BԂKW��ܳ/R�D,�ٌ�{w���ko������-���&��5%�bI]�4���hƅ;�%˺�	��{b:���~�+s�	� ���t�����C��}����,JN��o�m�����$2%͓�gy���Ĭ�`�QUkQ���drG���>�_��{,�Ȅ8�ʌ���ZS8k�%���%%�cde��5{����a�M�W��6���H�'�/UU�,ND�ˎ�Xc1ƥRf��x��]ξ�o?���[�,�lv�}ܶ����{�eh7��N���b��&r���K@&�ʔm�dB����q��1���|�!��S�o��{�S�<�g�c��˲�{���3k�K99��ǄV�u���>]�[#�2�&4M�F��h�h@KP�2������4��A����ѷ�2����D\$i�<�2�UИ��'��Պqs"��1eK�l_�m�$��u�\�b�2`d@�J�6�\
�p��*B<Fc�].8����s��]��T�b:	 ��sR:>��>9-9H�YV�)kN��m<��X�X�<�����&��J'k(�u]��[�˖��&/\��g^d���t:���f�C���Sn߾���>�����m�CX[P�wo}ć����6�x�%�ַ�|�
���8%�u��α�{���m���dv��{��[?{��{��G�!˦A���1��n�ܾ=���?z�g�~�ͭ��r���f�(+�i��|U�	���?uz{l]߼9{��b�:&�,�^�`���w���=�x�DE>���:8@0ƢQ��v��_E�R%�D���Ύ���~�'�Ϩ����vt8�gM�=k�;�^i0Rc�#"FL)��J͔eM�4+M�b�|DGa�Ŵ�8����""�(J.^�e2���ܺu���^R/	D���c�i�"��!�&su��pѯ�����2�=a��\[��s���#�1������ں�p������:)+&Q����س���0'GN'z�y�
���������h�ӕV�@J����ضH(\b����рyL�\)��M��[�a8�����'+��n��8�1 ��;e�Z8V�C
/+Mwo��Ꚏ*�7K��1�+�i*�7M�~�l6��n�[�PR/�(�sx�4MK���ǶAU���D�+���9��7_��o0�G�.��쀪�N��|�g�í�e*�ý�/�u��da����Cvv�S��b��(-�G<x�[4�&��WQ-9>�r���y�m�}�����K	56շ���CmQ0�����9�� �:A}��e�6*M�1�g�)lnm�s%��m��j�]��E�@?����@z��j��E�z�iA��2ٚ�c
��A5�i<�3�^��_�����[�mˤ2�P�Ĕ�g$`բ&�1P����s|��k׮��������p<_b���X�h��b�p��.�i����7�:GӇ��nP7��2�r�bI�m�lǷs>����xT[�-U��	��<9RSũ1W$�D/�G��yj�����y��7����!���:����>˷n�����~�мȄ����,%��x�����}k�rs|h՘I�X�{�������O��l��v.�{8(Km��
�p��ڐqU�Y�$�u֡eI)d��]�<�U��2Q��M�\��G+�(J��91����
��|�lv���>�	�BI�xM{��D��:\�J��9]�w2��t�MӜ���癥˝438ι�d��Nw�0s�n���}��u&��?���w>��x��d��Y���b[\QUɠ5qUFsU8Z��)��{̎7G���e6�i�}�w�������Z���Cb�b��Sɶ���~�V�6��9�H)�v ��K��=    IDAT�󂢌-U%XI�/�7��t������;<|pH�R�$6Ɉ�J7}:���Jr��pq4>�w���$�����`�h4�(�����Ո�0��T�w~���D۶�*�*��?{t�\��loo2W��o�펊���/��4�n��0;f6;b1��6e:we���;I��E�^(�c��=	��i�R�PI�
Ԓ3�U�O�7�O$QM�1��TU���:��,.��Р0�D�cQ�?#VI K��t��3��z�J
=��!�HE.	��ǧ�j�d�N���X�Q<�E4�8�H�^Z�5�%kEmm�$��j����t���ھ.�_1���]_4��4��c�z������L�X��;�(0��e2�P���EY��D�BB�T�W�bF�������k�w�F0��11��Q�D���F�Z�4���UgQ$�rY�U�ӦiXV	��m �S�0�k;R�i��׾��?���O:}���aDR1�ު(w³(�b�Aۦ�;;;lmmqtt�b�X�Ķm;�x����\E�{��Y?��V�
�e&�_�h�#��We��t~}��1�����1�q:��y���E7����ĉ��9�>������m�z�`9;bw{�A����s����{g���;;h���뀿[M^Ʉ|�Y���xc�y�Z�A���Bo`���r�<-���$c0�uK��>;:���!���L�3�`�vL4�95!�Y[1)�0� Q�<�xz��9�-0Q-�VT� ���E\ǔ��I�o�G~ͷ'���S�J6|��U)DS�w�UG���,t�p�V��(	�&�G�g"_�nO@�k�K�jQ,F\yS���ֽd��<݌@V��dEJt�
bH�;yIo
�����&�Fl�RFULt��$�M獧���g�@��1QM��Jʚκ�cҼ��P�t�"���,M���,@S���M ���q���5ޮGU��Ԭ�^`92c�5��n~����������"�ۧ���{#Glr���QըF뽯���u�ʐ��Ȣ��E�	��_��{���l��h��kj��%�+�����v,e-�25�%�cM��5���q�Ĺ%m�2_$/�A5�m��a8�
A5p�������H
��h�Ƞ�VN�3Eߟt�d�Y3`i����]nܸ����*���F���E~����_~���x�^Ɯ�M��h֍���5?i�R=�˸��g���iO�%j0�+�6��xk~ĝ�c2�ę��#�z��E�.��{{ܽ}���}Ignӵm�l��9W��k��m0�~N�6m۲\���6)S]�ǇH��mX֋�6��i��b!�[�,ʑ�M�H�,��(�/+�(!%�4
�8*�E:%z��6�3��$4���,yf�������мc<M޳�kڦI��8��J�� �rzA#^#�J���q�"Z̟�v�IF}��tL�t�F��
���n��u��Xm�+!�)�!/Z,��t/�x��K<��M�Ĕ++練}W��9���Mn�!��_����
�I�e@L�J$6(.�-&� �&�W:��*B�#`L��e��"]Vsx����[N���n��[�������ϓ���s]β��gK����)���0�/�1X�Iy�Q���c�Z��n��E�|�>f{|��L#VU��Ԃ4U�/A*��t2J�Z�B0�	>�"cbǊxr�+�sFՈ�p���)ꔭ�Lg�<����w���/pt����{��ݻO��:��N�/�Ϭ^�~�Y�,��B飣���N2�����ѩ��l���������s������ڧ~�3y"�p8d�X��˙A:I��x�ܕ��E��ΘNۗ�K!�\*ki5�8>`~t�C[a)� �6+0mM��ђ��Bʮ�!���٧��������LA�����m�jB\"&�
�u��䶟����Ҙ�#c�M���q�BL���R�T��K����4�,��X�5.U=),QS�L2>VK
�8Q:�����
N��Oq��º�C3�C����FYU����X��;�I��<�:�b�ˠ����}��
	jL-&`5M���N�������8�>�n��A�²��&+�&�E�H�`<I���\�P�3�M,�1մ��k�twh'l�E�I�ӗڸB��x���S�IxS�t����(�2(v�7џofVK�'KD냾�����Y������������r��Fl��}F����''�ϸn������*Re��,�ъ��x�4"̌m� �ۋ/BVߗ�c�'0}����j�O6�F�xYSv���F�R�
c|xR6�����e�hV����;;;���k��|�����&�	ՠd>����z�rѰ�l�8�V�&`U�,��Z,+�g�a>�����b���J��[���j 'U�4�c�`-gg@����,DO��;k@�"��~[�5��1i�������&�D�3����%�8l!�o!�
�@�HL��F�h1��L�E�4I�^�hh�TǖΔW*��^*�
E�S�$��İ�N����Θ��Y���ghi�b���,�N.�ze(��I�H,F�Nq�{�*u8Xy��{?�IY�Ic�!z��4�jK@ X�8���s1�b
�kH��D�X��[@�O��c�u�}&��l�2}��AC�}]���L{��r
�����jNd�;��a�3U�0E2�&U��@$1	$ÞH4i�ŷ�U�FD�">���b,���B��+�gH���;�]�ݑ���%1��0�C����I�Zs��Op��Aߺ�V��y��o��|ǘ��ׯǩk���~\����i�q���y��ַx*�3j���j�Xc�a�%\d��b���e�B�sA�tzE'�N��G�APO�����?��
VI�&�
]�\��c�cc#�lU���[o��o���\�t)�������������Y��(���T�N��*v<|�p�Y8Y�z�W���;d��3v�w�W�9�������'2g��Hh��h���Q����t��<��}���_����=�ɞ@m�]b�Jg!�2݌PR�Lh �� &`b��M�8am7%��b�w�o�k���_R�S
o�t��$�� I�
�J�4D�D�'��N�f|X"�슧��$���O�7&%�k*����Đ,[\WMG5%�� ��R=\���c�`�&�!�im���&��ݦ'T�vá!�F���\������`pj1e2ê�Đ�N�Q�m�����y��;o���k����U4'a���8�l]�Q���5�+�䟙A����S߰ޘ�?v�tw]��d�1�99^%%Y3�W�I [$+��eW
7{T��>g5,��[,�.�����9Gi�� �l� /�'����xw�+C,>+Ě�=u��`�ց�Y���y��B��\g,}g�c���+���`DUV8c�1VC�qv�"�p�h���wŪ�K���Q;�]�:��=E%���Ah�8#���t��-���v��y��:�`���dBU*GG3�ۻ�|�����Y,�Õ�i8��/r��e�����Ν;ܿ�}ˠ([f��t��2C���2c�����fh��B�n������g ��������=�!�b�l+�{�;�}ј>��][�+TU��]�P����6��EA-��o�-�2o�nM��dԢ>U��@��r5=�F��d�L
u:��&9ƈ+:v%�41R��#�׮�+�����	��~��VU�eC�6����/`�`]�(�.I:B��[ �`c��h}
����m��ʤ}5��>�QbL�/�`�+Ř&OԆб����;�I��bt���A'��+�>�?�yzb����*���#�rw������YgwO�k<m��+2�H�L�QQb�ћ�`�bR}��'�I���+ �IV+10'�;�poDc���KC�I��;O�|�������y5�巜��b��cy���g�}r<���g�_;+BsV�(��o}ΥJ5!x�5��c��	M�����7����:Ř�&�2)�������S���l��v.�����`&1�E0�F5�^�7���Ƙ�~���0��T3�<Bh}b%�j'�� t���hs��9f4����n�������&}t����՗~���[�xq����|���{�{ꕯ��dbT�|��+�NUW>Wg��+�]�;:���1��:r��#�����~ˬ�j2�uα������
�>n[���xU�7g��{�U��mR��xT<1Z����)�	��XpE ���`:;��E�	��]����g�V�ڝ�'�W�0�_�Aȓ�Y�K����d���pJ��Ԩ`I7�ѐ&�2�P#fD�w�ͥ-��UI��v�%b��u��<?�k�1��u����Y�_ak�E��t�DR �m�K�S���z�fxW�s���哄���bd�)7���@}�n��ۯT���-��6������^q��?IX���%v �v��4�$�r:�#���	gA�S�$�W�����L2���OK3�B�k��}���V�# �&��9,i0EEӂ1���@S3
���x��2��c��q3�2�7"C���K�_-�À-��Ō�[;4�R�kv'����fH45�)� Ô��˸�|��h�u����#��c��,��.N4�����$��˼�`��d��Ax�jk�p��.1�0��l�mB;$ĂڍY6J�~���­Ch:_)TlWkA�I�$1B�uZ�k��0� 堢�*|�Kf�}"�_�3g[٫/�Z��!�r�Hظ������]���ǝ
g$�B�S�Nk	�j
��q�H��4���E]����;\�t����������=�/�����s3�y�g����'�����v.���ى��)�߫�jEP�Jie���Z��:��F�;���3�-988�iF���!��>/�r���vvv)˂�tJ}����ի<���:�����c{{����GB�O
q�5�v,ow�����}��Y�3y^8W�;�ugc~��
f`��/g\gP�}���U�izN��az�?�cߏ=�!�I^��ʧ<���X
�)}�#�Y��[���Y�~���)���0L�9}?���HA�z
�Pز hK �k�C66��-8n����[���g,.\����|�%�ج@*�&�RT�;�`c�.�YR��;u����u�����\nQu�M=��=�/]WO���!ee�L�eX��;�0�K�zsG<s�;�Z�s/��rx��ͯ��W��
�+,�����~�[�7�~`o_��,��a�F8��J�X ����嫴m���{\�v��}����w|�W���Wee�����@#
[h1qf�x��ח���}����޸q#�m�y��"� RkJ���j	�Ɵ��q��t��2w^�	�3�p||̃���u�dr��G����?���o������.�����Y�7����ڒ�(�r�J�]FȜ���AOX�Eǯ���?p��?�K:��b�&�����	wbS��?z�EO�B�߳b8�4(<�~�-��-�b�2�z&�K�^�������|+u��3e�ѝ�~XىH*��=�V3]U��kҎN��S���i��o]�q�ϟ��ڢ#	�Y%���$��n�,V�,�Q���zl9fs��q���!���H���%֕X;���H`<��5�˲iPM����Г,�Q���%���P�����"4U�1����s�uU+X�5���Z���5��%�	��)�%A5���#�0/'�Q^�k�>%Jb���'2����_�>���l$��_�i�@-�������K����?]��ܿ9Y�w6Mr��
<>$������D,��ߥ������7�����d2����?���q|<�M��EӴeYVQ���HlU�i[��b{���e�B��f�n,74�&��H[�i)2G�RU[M��QU��VTN�T���:����ASČ�Ѫ�fs��e��px���k��s��U9fP�����N�ݻǝ;w�L&\�|y�ӛN��t�>K�;t������ߏ�v���e��������}��{���_�c��S@����ǲggl��j}���Q��S!���>}-c��O�2I�g��u��|҈����Gx���u���y��9�><���Re��>(����@��{��k���>���a�/:�%��D��/����S�K�� e�ŕ�np��5����̨�c���S�o]�JA3]2Y���_����M�B��*��O-z��uD1x�D
p�M�Z��hLY�ƭ�_�釣f��	3���@�E�Lb���'[1�k�@�!�-�Iv�j�	,j��骫��-�O�����\�u�����Z\���~��>@̥<�����=�#V�QJ�����ژ�)۵L��Q��)�[�<���/\��'���w�r6��?�F�F����g���x��F�>�H�=
?���ѧ+��e�\�sA���������E�:�u!%nȑ��*^U�*ASC:C�U�w\�L�ٳ.�RX̑+z�z2r��-<x���6��&��pLQ�)}�����u��i9��[o�|���z���:��g�2�9��Fn��C#9�7�����~bM^M�e���+�Ē��	[�uF\�7V�I��=������$�������r'ӌ����g9�kǄ���:)������}Z��^D#���]Z���Q}K[/y�͟���S�˘a�`p���ã��ܾ���87dkwL�i��-�������z�Kw��!������wߡnTO<��GZ�u#�@aS8�,u��:eoc@R&��l�O��1�_;C��5��B��s0E�+�P�T�ͤ�Wlh0aLԐ�=1Dծ�!����h��2�N��9ۍ��>�g��_�������Ҝ�ѷnY�w�y����Ǔc:�8{�����n�m�(+bT�&�o����ʵ�?�\�����H}�\��nx�޽�nw�b[��C���zUDE<Q�3eq��|��l�������_��M�֭[�+���\}�@����s( ��X�u��ߏ/����֭[���y����:��DD��?��qm�M�����j��F�eT���P��,����h��S�C�D-֔�XB�GC����������
�;W�پĻ�!����)}`��p8<�1�����H�|>˗�� �Y����ڼ�q���g���Z�h�rD�g�����w<-⪪��+�׿&�0��^*��=f)�(�~�TI��\������|�Ӯ��J�;���߫��||$�˓��'�\��˳&�_�w��67-Plʎ]},US����o�����h��k�|q¥���R�Qmy�����!�1�ł��+|����W����x�*�shU�\.�O?�?�ɏiB��
TQ">*MT�
;�nCD�g-Zv�%��Rv�*���m[�!/^d{{���ͭ{�C��� !�H*|]PT#�	�(Y�|hS�{R�$�HO;7�L&���7(˒�tʻ������^i���c_�@__j����c�ia݄߯�;�{�f�8��eM��,K~�6�ؓ��k�4�C~���L�\��'�p?�?8�z��O_ڽ�Еû�ãoq�������j��h�r����[���h�Ϭݼy�ܺu��n���op��ݹuK�_��@�y�62����U�P_���o~��͛E�M�`n޼�_}�U{�?������~n޼i�� ������z�Bw�N/\������E�p�:���������Z������GGGᥗ^
���w�<�����h���=�;1s�F�CsT�&����#�:�(�ӝiW1ã*X���\��y�7�/�گ��y���b�Ac�2/��-�����{R{�w��Px�wvFf���5g�<x�ߵ���qL�)���`���$\*g��_t��y+P�\.QMY���'��V�	����S���~���7��-�� ��#�r�9�ڱ)�I?`�Y1ۻf����2G_��2w>�
�/��ϻ�?��!��W{Xm�g����N��bwW�    IDAT4�����#�#�[�O1(6�r��(����;���䭷ޢY(UUp�+7��K�o��l����H��1}x��������oػ� �A ��5���BU�o_��Oږ��i��!��t��6b�ٚln������K/q��U�����kNk���h�����l��:L�lm]��s_g��s����ǀ�M,�I�ڳ'��W�~�:/����ܺ�Ç�<|��Tbŧm}��^�2��斫>��]x���ni���]���Z��p����e�z
�|�"O?�����)�W�v.����u��ۣ���xn6�Q�����L�b�+e��Ԉs�w6P�!L�o�����oKR0����s�)�[G
��`�;qoq���u�������9Y�	M�������^{I ^~�u��n��@���\}�+����Ķ�9޺  ��L���y� 	����tl�) �	5Ќ���rA�����a	j�_w�E#/����͛���~�e�������a�ؿ��! �H|(�O��ݺ��2ڑa�?*b�{��{�˲�"��Ht�;Ｃ�������Q�����*�(��XЗm[ԧ��"RG�V���q5	�����V�ie����{�:	�@c�唷�~���S��;���[��S��s1�#��h%�=ku��t<쭷?Zg��]}֭�ֿ���yL��1�u\^��_�X�����e��gn_{6g�>�=)@���p�դKD4yΉb���c"��H�!gN>��i&]b��~�_��3}�x@��:���{�G>z:�:�/�b�̧kc��ܹ��]�Ե�\�x��4lo�p�ZIQ9666Mvy��wU��o�5~�����+ϲ�<�ǲ�y�����������}���6�MR����Mb�)�Ոrc�_�֯����o���t�ҕUJ�e5dkk7��+��7 �@m����ä�>�|���]��$F��f1]�8^��������o�w�"|���⒢H �(
&�	���\�t�o��5~�~�?��0������>n>��>�̶]}��`�<�:�1��<+�t^;}_w��c@4U�bS�GUÊ�W�����ln�|$���უm�}�k�ݿ����n򢭎�iƣ����LhC�3�R]e�b�����=�'���?��!$���͛�$z~FK���^{�%y����֭kr��m���y/ ��Ƽ��X.2fr<��ӳ�����/����D_~�o2�V�.����`�z^/���E]U	��K��+��m�r�	UY��~$US�c$ �F�	CY��m!�h����y�^T��j��ea$V���R�S6�����Z놮D����V���6ŊB)��.RH�"Έ�a��Ęo�����b�ۑ�'������'���B�Z;zX�U�����w���p��M��},���ى͝&�u,�SU�ѫq� j�i�v�VVˢ�Nb*��M�u]�4~e2�+g@�6�L�]' bp�ć��Q�;��|�`g�2/��Uvw�y��w1����,w������u�v���s�}�m��Ϯ�;�\U�{�r�\���5�����e}[Q$ֳm�UH83b1��NF�`�;N�
ׁ�,`N,ʲ<��}�����{�o_�G�1����Ζ�@�7bp�2���FTU�tz��d�]��K�1����*��E��
cW��'"kш5��#��ćh��I�v�-���A}�hR��q��x߅�K��&����Or͞t}�lE������-"�!����bڞ������-t>	�[�3��;�N��s'>�"�����.Z�3�#�{o�.���=�ۿ��F�S�����n<��zIeGLƻ8�}H3S�7�����������3��S�uq�+*�Ұ��.��?�{̷�_|���A��k_�j0fk�����0XW�\IQ���^���*���7ٹ��r�d>�a������w��.���7�b��Ʒ�O_c:m�ؾ�׿Qp��g���}�>����C*�E�
����|�2[[[�E�1p8=��*�޽�|����vY�ZV�zHz"��L@���u]3�1�HF�ѩHD#�}z=���#��xU-*'�d�轧��GBh1&eE���`�*bPE:�m�0���~1�l>}�ҥK����O�H��������ϗ�[�������m1jcۺi6
W��Ъ��^����v����տ3�b�x��A������W����#�o���@ �������ZJU��V�TE-m��Jdo[vؚ�u^���G�~;��33�@G�)�V�h�������j�6�+�_�儉�M�)CJ��z�CE��h�X34"v�Ī�¨1�Ɏ1&��� �1��Hcw��UF�h�NJ)��F�T�7Vŕ��B�
����/��FS1B�9QI��(�b.����c�U��{�1��J�$��9KԈj"��%�?>|��;��f0(k���]1o�{�e�����"��q����UUm�����><��������$�I�[BC�Ӂ>�^��v~mXn�@c�m�aU�@V�x�z�]g�B����|���ĸĺ���>��./�E�r�h4�|��+'4џ�2HȃK�Ԝ�zM�>y�/Z�����BL!#��d�cS��XGaEY��mp�`�T<=�7]	��q&�+�D�U$U�ǈ���U�j�&��Ŋ������CK��}g,���kJ�݂��l
s�Ɣ)fU�U>3���o�"��b�w ��j��ekg�2��$@2��Z��cm�u��^��Oh�oN_������u%��h v,r��p�w���w�������T�
��&4QM��p��S1,+ں�駟fcc�b����|�������m=�G�6�2�Lx��g���a�\�\Ԉ�ˆ����~�����m��Q�>���{�R��_cwg���-�����6�����W��K�N�-'c[�-���9��o�����'��5=�ym��}4�����0�%8���m������?3��W���̋Yc��g
���ǖ�%�,Q�:���Y̗�8t�����n�_�n�AU��h4x� �/^ؖ��-�ҍ��[ΚƔ�T��Q���F5�\�/Ն�YiŗfWd1Y.mٌb#��P|S�2nצ�%���cql�غ��3��`�C#3��c�##�����DA�v �T��0��m����hCB,�ja��0*Dba��P)*ވ��6D�J��3��łE,�(�k�Q��M*Uh�b��(xm1Q�xL4��8)�-�q=�D�U^	�Z�$��hX�c79t��=Fl7����|"Q�JFa2i�ȉ��b:���Xi�t�T��,T�:���Z��ֺ�lCx�����^�ڷW������WL�K��R׷�����~�;�	��ED��{���klZ�N�6ޕ��|�Wn��҄`���?ab<�1����?�hW�ҦbھMu>�*!�T���o����~���;�ۧ@�����3,���>��0�:�x۰�r\7�NV'�Z�? �͠���
����_Ɩ4q�B���U��� �2���d��d4���%�ii��K�6̎���b{k�j8 ����V��ʌ�l�(�#6-!$?���p� kS��������ɴY#8gp��XF)�W����s��G̎8:�&�Zr�zM��ve�>�a�g���ON���>���?�<������Z�=�qw�C�F#��qVY�,x�`��~��s<��|��lmn ��m�x��2�s��}��?����G?��G0��(����cBL&��P_Ӵ5w>�,����W���^bs��h�W�C����#�{Ɠ	M��=>��V�������;n�y@�JWR���ʲ]�`���ɐg��A5|��xBi�Q�BY���W���z��\T�9ӣ#�}�O�ٛʭ[�0ư1w���	�13��9��#(�儹�������G�����l�Lp�b5⌤JJQS�@��h@�*<���(���h�����bkk���.5bE�h2���(�����-�_�H�ث҆�mf�/�Rc��f�����Q5����8�1�oC4Xi%X+�x6��v�q�k[� ��5
�p���'�W#XREK���FBT�i	�k�cpEAT]�1�h�����)�����1���1��dzL>[ɲ(
����MB�iN��(���H�(�����<���x@�%eʧ�4���S���7��z~,�%��9,�n��e|�ò�:a�h��l*-L�Q�vP���I�K��Z�����z�1�V�ê�6�Ν;<��4��W��\�uӨ���=����,��* P���	8	��X
��Т�Q/g �*b�6��T轡��?}�M���ݹĥK0����/�ı>������Y���9�Ұd�q������3}����`��Ƣb��l��8S�6��W�����p��.�I�d8��-A-�i���m�߽�dk��y����y�L��I�;5)�k
Ga,�+hb���X��eQ`]*AU�m��&c2�1� gk����7��$���>g��{o�YYUY�7�E��Q�Ƃ4��@���������E�e =Λa@�0�a��戶�#Q$5����ޫ�����.����q�fV5�ZlJM�Hd޼Kč8���~߅v>���y��[���}R�H���Cj����Ϻ]���ϧ�>k�����c���p�Z�72�u$�X�����֏���c���Wv'$o��C�p��G����-��7����+Wv0�,}��R�m�K�����-G���4-J�O�_�am�)ʂ#]��t��PJ���q/�b	>���������>MQ�� �cL�-����}f�1�g��S�y|� �uG���Jcl��N�|t�.���w���b�]��R�Ӑ��R��/'��X~ު%�Oz�R��,P��5����L���>|�xTR%ZChm�$���,)^|�y��^�g���}k5"
���c��'''j6�G�Ь���!xΦg�m��S4vL�>4"1�I"��Y�8��ql��P���F��Ry�4)��Z&�Y�I	b�q�齂5Z[�Ŝ!�k����b)e8���^�1I��L��
�"Ď�d�QS��&��cDooF���~�1�R����-_C��J��q山*c����,ӧ,)�?/R�$	��N֪�bAb1O����w������|>�(���q��5��L$v�m=�RZ��{��ۇ{׮�ͺ���Փ���*����S��[���~���KӅ�c쒮�Wj�B��4&��Rk����#�e'�%�sw���$�a�i���}���4H�n������h������2[�ns�ib5���>&�|9�S*[�el���i2mC��I�����dl�}��aP�p�7��˽ֱc��_�_~���]�a�V2�J���ڶ5,�sl�c&��{�y~��W����l�R�y���~}pW��5Xm�YJW%�B�ǐ�g��aB���8g|$dQ�����kLF���~�Ǆ�e\!� �V���$���Q�iړ�u_�>��.�o�U�Fಜ�z٠�ؔT�АT��<Ea��-'�;4��t�l����?z��+���r��{��o�?�/�e\e��{��)�fOX!�.�ܑ����]�����]��\�5�_�썶�F%���:3}C���pŘ���[o�g����{� �|�J��y�Z����)�t�����%��]gsm�����h����,jR
4������~��?���Kl�<v�O;.ϯ���mۢ�����rQ�K��sy|�s���{>{��A_�R��g,�9��o��W^��g�ak}�_|���66��>���C����͙˔.��E$,�?�E�0;;e��7S0�L@ �@m۲����%Qʠ�,��Ƹ�{6nY�L) 1� ���t�A��kT0�0T줘mHR�������A�)k@�����rp��2lF;��,�gȃ
B�������(M�l$�\*5��5]�0$��2dKt��yã�]�o�s�=W,�;�FS6O�èIHʙꔲ:I>~ou�7�DT)�W�@"=!�tm��	Nk�LֈX�"��+���>��i$v��cR�h�"�d��y�~
PΟ���Z�f:�L���l�b$�K�D�T2�U�2�s���灐�b3�q�Z���l=�=��ؕEŃy�G��r���X߀Ã'3�(��U�����=8s|Ri�ݡ4�*+�XIL�@m�ȡΟRPy^jX����Ӷ�c�D�(M�\:��a݈�_�%����x��g)�����SG���7�r��u�z����{x��S\f�����Z)S8�����=
ED�mA"���\��~�|�����o�)0v���-^y���%�D�,z�]��	�$$��3l[[[@&E5M��p\�,��� ?����������MI`�j�DD��"���[�u�l������c~�_�����IL*�IM�g\�o�X���e,�AE!rvẋ�}��]q��1ׯ�0����U���m9;;�YM����;��֛|��m���ZML9�D�
�I�tDbJ�2�[�ܻ��ݫ�nl�QtmK0��D
M�/<z�����cP���5-���m�t���@oU�XfE2p`K�ד2}����c�����o8ހwW2em��ս�vm�/�U~���ʋ/=��x�o�I1��r��=�ܻ�b�@k(]%9��B�U��$m�b���6@@���uH�h�~�$�L`L�<��>�ڈ&�{v.E�ҽ��ܨ%��h��!F ��V3�0;�^�NK�z�(aI�QY�{Ũ@kM��sMU�Y��UI�JΦ� *�K;���ͥWb��A`J�y��HKJ$���%��m���zi.��/�����BΚ&�
D�Z��lS�\�>Hv-�]��9��$�m(J�-T0�E��Vִ֕�n��!Z{"U�M?x����x��:��e�ү����Ԡ��͛�����b�C	�AL\H�_��!�����hKf��eP103�Tbvn�j��c:�Ҷ-���d?ĵ���O����k~�7�ĵkW���:�0 �(���%�U��<Y�>ڶ�m�eve�֨4���	�O��}R�OD~^��}f���$��߱�q%/��2�<�[tM�qt�iy��*�:�X���:89��)1�H�cz���`M")A�6e&�]T���c�ꀖ<Y�$�63s��1vFU��`L�}T�5���(]v$899�n*���&�?�V�K��GW]e>�������-��Kr�R;2�~����w�XD����K��`lD�fѴܾ9;����Ӈ<��#���8;��RYJD;K�36�Y����	�*)\)pvz̷��/X[[cT� ��>�)M�55)vLώ89="����x7�=�_�P�Đ��$�ȁT�8�rx|���w(]�����W ��wl���,s���>����$8mxZ�Հo��2(*(����kVE�/��e��tP���X
+E���&�W���˯���̋/����6�-9;;���qp����I���5&eE�,��@d<Z��J�F2.�g�Z��k�L�3�z��#J��l��[�M	�Ǣ��2c�Gi��*^)d̲��#,�g�L>OԋŅ@{(���R"�\�,sŒ�R�ݘ^�h��J�Ϥ���y��R��#�@�ۜY����;��R��,9�Н�\�09x�1,�K��u&� ����H�
LH=�C+��ω,-�͘��H�A���%���)�K�9��DY:�Q�Zg��h*v��	=
^TJ����>|xT��u�vۊF���*�u�֧}}g�!��إ&�i܅�3]�"�EU��}��2�މv9Xr����g���2u]g*�����Ψ�*�y����`cc����S���vy�X�s|R�d�<,�]�-%^Vu�T�da�ՠo��w�?ia�y(�B�陼�īuΪ�!E���v-ڕ����i��,������ѣ.�r�
]�]ؠ�uM�4� <�b��{������*V	��k9����*7�^ac\H4!g1|��NV��*"@� ����~�V�����������}�ٽ/b[�Vk�*9���В��[X<M�,    IDATsF��8�8:9������\����t���+	���f(m�L&�D���Vk�V9!�-��&�LP=�H��ZZ�*JRt��Ih#8F;B�X#9Ќ�A:0d z�$��>�(�)�����k[LPH�>h�{�M�u]c�f\U,���tX������2�N�J�����q��K�����R�i�6��s٦����g�ʾ\��\�C�h4b�^x��ۿ����Z>��>��0����՚�|���!ggg��_�%B�fQ�PJQ�%�;�=�2�s���>�	fYB�{�lV�]&]��(3��țݔ�L6��~c��>�U<k�D2FDHBO��k���s�/%���(T�	1�e����k=D����
�!�#��uuX��\-��1��91$߷�D|.�O���,��]:�Pʀ���S����fx�����x<^�������8 O0���!�{҇��@� an�B�����6ڇq]�ηm1_̪���ַ�_�㣟_�*��~�c��F�I��!�����cӎ��*A�.�S�똢B�`�M$��Bk�B���g��ʸ������.N�q��w1�G��2�89��sݱ������w��z��2��W��g&�	Mӡ�FG��:/�� 채�>�*�y���I���}Q,x�)�H�<�&�e1Bk�'�>0��:|�ΒR�M� ,�g�pq=�M�1�@Ȼ.���b�DT>y���Jڮ��c�J��H��q�1d��s�%�y����/�)���Oh�\�$?�{*�	���3l�bʒ�K4~����OL۠;ێzq��?x�޿���X�1�ٌ�b���,�3��poL� $O)�Γ�q}prF�����f�`R�"����R���0�Цb����^y�����^f<���#f������c�+0�X�P��Ԣ�`��k�$����-	�Ǩ�C�$�ypvL�E�WH��)���s4O�߫Y�լ����l (�X5��Hm�H�s��P:au���)��d ���\���Y��:��u���ɪ y@e����'_�Oi.�����Y@2��.n�FG+/���� ��~�dܿ0�TU@K��[�������5B?R�c�B�R ��M����W�,����{����Q��>���������Q_:,������Xl��q���{��f��L<�nnKt�IEI���Ǚ+-h)ʼ�w]ۗ\=�����lpzz�3�).���L�6���ec�2C>l�677���㥗^�W^a�ǜ||����CX���98Q�tI��ͥJSN0�-�1��Z�����欪*Du����r#�Y.����pơ�b��
EL�D�wC�pe�[��)&u�q��K��&0CP��h��%��r��N[�3'!O�S��F*��O����=ñ�y����uJ	����r$��$GW?ؤI�8�|��1�D���i��}�����ID�d{�e���$��j�\yC@ň��|�R҅V�`��U�k3�ו�pvz�N��֞NO��3ƚ�Y�g�y��=�'-�Jb�����Q�S}7o�L7o�q�ԋ��AI=�L�!	>D)G���$�8;��오 %�C�	H�����䄔�E͇wnspp�h4��8<:�J)��)u[c�S�~�m�����3�<�̦���1��!S��]x�J���jľ�.�a��ߗ變���!ڶe��.'�Ld�����i��6����Bz�=vy�_���b_��[�@�<��rP�:��@��.ι~�]>�{�G|������g>] �6��4�C%A;Ka,I11oj�6(k�AR�@��i&��gM���&v�7���T��d�aM�i��zA�,�E��(2�ue������Zj��&���������o���D�2c�$��z����R�$�p��h�$��gQQ��(ML�#���XC1Ҙh3x\G��^J!KH��AZd�hⱅaTd1���������)un�vy~��۶���ev�m����M���Ӵ�VU���ll��t:�����9��������UU1���2�N���9�������9���@Y�,[N���H/�;��$�C+�1M�\�T�5���!B*M�µQ*c�SPK��2�ѯm������,^9Ɠ�<{Ѵ` Y�b I��H���W��(�Z-�'�$b8ߘj�2�^�4EAY��ev�ϡ�+X�,�f��H�xR���������D�QHt�H�.�XIT�c��pI"�:�$&�5�P.��M������"�����J�$ҹ��l{29�R�#J�[��O�yL]gT��k/�S����w��(�V|S��1�&��t�]B��ipe)1&e�5�+2�8�Z�v���$@
W *���I֧�֖ʍ�WUf���(��o�������}�Y������1fyc����KA�%-�U��0ПTz~��-�N���?��؞Y�rY.w�s��A�H.�̯�S��L������3��"�i��\��dw�����9>�������T� a������os|4�t�;�����A�+U�Y�͢fT�\3�k2+�B��tG�����A��L�ߚ� )0��Ѩd2{Weצ}���C�/K�1��.w��)�jV��ṡ=}�XeI�u9�c�J�.�B�&I��8kp���U~l,�p�a��jC<�u�"^Z�}X�v>g���j��	j��E�l���A,ZU1��Ç�<�LC��UÆ��nX�{X�>�~���i�~��KU�O
���Cw</m /�_��|��5�ס|<ظu]���׷7��Tw�&W����&M�pxr�$R����3��E��mhЩn�&H@�E�yO*�ULA^�R8OzĔ(�k��Q)bL(ՓP�!��+Eˊ�P����}�ߺ��A�֚�u9�3�a��ƈR�IU]���ka^g����>j֞a��r=��X[,��(���\��g��\�UP���(P:o���m�d$%�E`:�+�-F㔱>�wI"��PS��Ux���N��Y�1Z�L�ԑ��Q�BJ���4����8c�c���AQUGhӖV����%^�w�o׋B��>�%��hL|ԺU��wQ��s������w�?zp��Ͽʯ��o1�w�fZ�I%Q"����.0.
�Γ��gKfuM)��x�h4BiǼi�ǜ�f��_���)W�^�C�tX�2�vri������3}���Cv�I��1���l��/(�vZ�#(�9��~�kb̯�:I��)u]/�1�=���ǘf�%����K�x��jИ��^��������&��[���g-��Z���K�so��]We�����9��BYE�	c���	�g� �b�T����U�� ���F��>upp�|:є�q��с�DY[ۦ���Jn�f۽m���U��O�\���KV�gi&���� ��v66؜\gws����̆���}Y�˟aR_��2*�Dl��i�(�
�
RR�ń���L�
5Ei�!��g�[�vX]������{�?⭷�����dz{�4d��11��$,�?��w���\�/��Ļ�T�6�K՜���0����d�����bY^�_��<�y�2��:㇇
� ���0�/�����z��l�9����|~ڟgp�4I:�Wh�PJch��}3� _�����:��F�eY�)8�L笣g�d��2�A�F����g��� )S$a��$�r�f�-�%8Pl��QYĺig�^҅�PBt��b����F��8|����eц�ۈh��s	9j��eU5��<r�RI�F"��)��ژ�� $k�Kb�(ZDy�@C��AsY��A:��� !�4e�C�uRZ5��F?&Q *����t�Gڮ��,�WZO��b�>��?9>Y�����uk2�|tvv�nݺ��������o|#Z�tA�mT��:ejچv��Ç|�{�t��ʫ_E����5zM¡mB�'��l~F�8g�eMΜ ���{��Xf���&J)n߾͇~����:��e�(1�zͥ 	gt�>擤/��S����o���v�)KCJ��K�=�G�L�ǘ�a�{"�Tp�s�]�y�
/��I��j[�S��˙B�;��h���N���1>Y���T����J	Lv�2���+3OR�j�h4b>]d����&�H[wh���V�R��O��:66��~�W�\��m�J�A�Z�lIQ�K��#?��yd�(����]�|:#t�|�����*D�Y ��(�}>�W�y�2T�o���W��	:o������.���U~��x��u�no���Q�rR_��iU�a�,��/7��F(m���^�'�6�����A��e�ch���܋/PM*O�xx�0c1����z�]�k�r��t��_���փ�k�Xt��@�B�y����[Y��*���`p�?�[x��o����:�Z��1�u��Ou��lvJ�4KG��k������nBX�Ƙ�n��huf5��:�?SBʏ��X�eV|r�tV/��j�`�!f۽\I�Rk"BL:����%9��1\3Q8+h��&��ߡ$W(4]3mU	Y1YD+���0�(�E��*�yH!%���䌨:�&���耊1�d�$��1��Je�B�Ť6�W���c�7�R�Q�R?�H��� ")v1�n4��z�4I$ň�DItZ���Q�F���gWRRJ�N9R�)�@�:��EQ�RJ�`��6`���F1���c!Y���=|l�����R,�v][We�������#�M��������NO�)���͛	mۦ(ʏM<⵱�j���x||h�|�Mv��g����]��DaQ�����ʢ�����|��tF�����(f����e�w�L�X,|����w�_���q!K�m��檧��Rͽ��0{x4-���'v=��cT?��ˌ������w�mH�L���������K\��1/�D��'�<�W�.�Q.g
����Z^�y{��Y��N_q���1�Q=z���&k#�ɓmU�h����d'�p�j4bwg���M���I1b�e{k�kׯsew7{��`|��{i�~F���ǿ�5=z�3�6�еs�����C�y�������>�ڞߣ%�xe�	)���|�?��b� ���3}	MJ�-*����+_�*���*���6��u7$\,���q��φ�M1�2�"�{HP7�B�P~��ӏ���@��w�;Ϛ���=�}�y��w���RYn�e�>��>�|?G0��U��g��n.��9��Ԭ�hV�g�˺��dyNC�ou޽,[�j��Im�����ܝ5/݅���������_���)C}:NNN�������l�����X�0Z���Y���|���6%"!%��m��`��$%ڈ��5L2F%AG笏	�V��*{�)QP-� ���Et�f�����[��$*DD�GR��9E�,E�����:�R-�)Af�譈?NAG�t��L
!:e;�z�/Ԧ��h�{�:01F�I@2�e�Jr��Z�C,�1��ڤ�s1�co�E
��>����AW�R�q�I:oA�l�K2��Ҵ�b1��8U��Fb�֒��|�:b8DB�	�ċ�6�I*��T$�BE��`SLN}*��[��	":F��Rڥ�x\� �t��!��HL2���M�
��Sw�y������w��6��|��.����.�m��|h�G&���j��*�M��|t�6��o�M�s/|���7pE��]h�� ��X���1�o���Gw	ƕ�MM�;�r��ƣ��w��?������׹u�V�yBJ�΢�.�!�C���K$g&��T��x��d��^\�.���Up�jau��9�d0�l.w�������W'�U��LG���]�Ւ>N�>wFY�N�>S���/�X���rPk2Á�#m]s���x�}�]�P=�E�ޕ�dbFR0*J6��xv��n쳳�E<"���2��I/oQ��^��!@%�U\�v���u
��8���7x����[ob]����V���=���f4������c��Q�K�~��xOkB���#�׷��ڥ(3S�	-�"����Ĥ�*���9�yՒqh�Pt�'&ͨ1M��UD��ʡ�%r����MP��Y��)K����mP��t$��-�t�� �3<����'a�T�!����WH�l�;��Zz����������w��t�z�u�����r�
���<��KH�q�����ѣGܿ���q�-���$�]�-�"aHQ0�����^}6h!6�	��]�6�4���?-���v�)tSRH�ke��Ց4Ac�$ʞ�������"�nH�KI�Z�H����`;���`;��N����L�T�E<�v�B�Z��C����͛7;��7o����������YF3�R�r�L�Ke��t�m�Z���}-B�)�I��6Q�eT2R*�]J�������_��$c��H4��N��N�C��%%��(����T���1XM, M2�A)���D�26D	$/1��$m�^Bx��,=�����VX�'�R�(U)cJ��	�^D��C�����(�]�`'6�-@��zܾ��k�֭[�d2�����3}G����6v�S��o$ԕ�	�4m[�빤������������7��ۿ�;���L��P"XWr��>���ͭ[���{[R6���zu����$�s|�]�r���-r�>��7}��;�Y�~�����|C�u�f3���@�x�JXH��f��]N(�I��30}VŘ��1����񒲿X,��j��
�]=��.����0�(Q�}1�r��c�Zf����s�RFH(��җ0�����6�@�iY�0��[��g��W��E��#���l�<VVWJ-˙Z.�U����^�!0�1�
$v�l��W�L5��|����>�U�{'���ccc���X�M�_.�>1���-3n}C���w��7�蒔�.%*m)ʒ��9M�,eo��ˀ�+�,)1�ϗ:��"c�����ym�����F�|^x>f6�q:=#�fm}���/pew��x��rL�\JʘMG�.�*c�zŇ���/���6Ta�F�
�x���Pn,ن�v �V\>k%d��֋Ռ_J��O�I/��h���s���>�^�h�y�l~��"�*
Wa�Ba(&%����`}�J}�O���ƍ�!&�x��G��sաq������x�"g)t-:"�4��3��d�>�L i�L
t
AGҺ�`Bd+A����I	�(I��1�h|��jQ>h���n��u1.?H]���k�(#���o�{���{?=��o�M;��IXخ1�ģ��Ye۶momS��OZ�N�k����h�8��W�0A�^��A���(���l�>�N���D�2�����$��BҺ��!im,ؔ�7J�����	ګ:�dt��+���""��:"��d�j�H�jD�����dc=��1�%�-7���a����0����<�G��>����۶���h#���;j6�����GGGR������|����g�͛7���3}��ݓ��BPb��]l�J����b���,f���G�l~Ʒ����s�/��2/��_��Wi������_~������t�h��u%m�b$��'�����#&�k4u�n?��_������]<x���d�`:�����l6G�Q5���O��Z>0=U<��[,�e�b�^<	�
�&bub(˒�|����d�s���A�o8�����R�X��놅�9G�$٢��	i����%��i�[c�f�R�=(��m�msV�y�-��tߧ�WK�O��i��ӊ�|�5��|�<�sד�k�
��8g�b�ʒ���Zm��l�0�,�:fӆ{\�,���(HQ�7-՚�Yٽ~b�(
�
�vL��''��*~����u&�1g�9��#�lsT7�u5���=��v�$�,	m̦�*�G�N���V��C����e;D��"!$f���`s{��G��;x�w�}���m�4UU�������b����a!lb��Y�k�5���3{:y��9=;�l6���
�_���wx��W����_Ѕ����[lo��}�m<�zE�hpnDJR@T��������S����.�~��=F����2v�r��c�\��kw�A�]n��q�u�1��ʰQY,�ι�Fί��z�j����������3�O(�x����׾�˯�o�q�۷?���^0����sm��    IDAT��Õ5�*{�lf������Y���U���xD�^�a4YG%�(�����t*v�(U8�.�+��קg���zWD�[ԋ��h�����uR��E�I	-J�I��:�3��%CM��E"mЁS�T��̕R��:��i�ME����	�ES�H�֝E[�u�Q:c��C�����d�>�w��ƍ��t ���tW�Wڣ��SE�(ڮR�.��Sl�N��F�I��騬�$�7:��ѕe�&���]���@Yy��EQ(����Z�ԳL&�|�?����1��R:�=R���c[��h�(^=�1e[����.�2�m�˿.���՗�y-�z���y�f��?��{��{I)�I��^�"���o��7oݼyS_�~]'�nݒ��뢔:�_�D��g
�nܸ!'''҅YD���6F-�Hl}}ipP�Řӳc~��-=zȽ�w��	���r<��v	�C����� ������g8UKf`�u��o�{�23��/C��U����Ռӻ�1 ᓹ0����m�Ռ�j���`�z;�2�0��`��kX����g���y��rPt�=��)�l�_f�rИ����8������m-:���rlݓXW�9��FL&Fe�f�_�LҮR�eT���Ễ�Z����Y�(���p#p���!��5�D�Q^~�+���qmo'��R��jD�\^�,����Υ���*����瓼J}ILe�Ӱ�J�
�\A�f3�Óc�z�-�����0�N�ЃA����,��Z�2�K�
?ϙS�h���"u3�mj�7�4�C�tݜ�4G'3NN�\����~YS����[;lnoѶ_�%���i2�{P��E��T&(��ڹ�PyY-��*\�/�jyx��q��Bsf�Y�c�7�{{{���s��RJ����0���e��5�}�Y67�������N3=�sp���GG�����M�)���r��m:�2��u�s)�(�N�ֺA̩��$/]D�7m7&�p>��a�����]���C�d:%�XGm�B֊�l������(������H��;���1&km�˔�6fjִf2��Η� �@g��Y�gG7n�P����������ɭ�o��o~]�c��y-���O����h����qP����p�{o�븷�'��$����w��ٸ���' �׮��\����]������g��6����n"J)�7�P���������͛7?���)�X,���RlD'%)���(���$�o�D��}ĝ���޻o�������8�k��Qe�ۚE�bBi���v.?Q&g���
���{w�����RD[CL1냹jI�0.{��<!�A��qy�_� ��eЗ�;�hm�'�:R�e9�^�����~�iJ	���P����.g!WI*���I�ße[e���U �OlI=����+�(H0��'y���Y/��'��y���]}���V_Z�,�٢��8WR�2k�T�ƣ5l��7��D1�1QY��l]�!�^�[����9>��Y	���H)��_��:��rA�S�.����1]����J���~�o��ݻ?�������V�uF�k�;�`�B�\��|����<�Α��iO1�a�1(�����^f:��d��o0�����C9�I�h���E��mO�k��0�\� �ɛ)�Կ,�b��[�E]%nmu��Z�}��.��������[UU���q��5ڶ�?�w>� c�Q�+ƌ�&��g�n��3���w�srv���U���_���g���Z2���G���T�k��{�#��]�1��^z1��W>%E���
>mt!mn͛��jT�%��֣���6<x�+��N�y��jp�IT�Ϸ�op��?�� �������F׫�t}U�8;;���}�5d�>Y �)��g?�����7�xC2�J$��Q֤�bL�ֽ�M���1*K�QI�����p����[뛘�Q�����9;�*�0��l��*�NO	OY�Q�}̥7��!P���|��P�a���<z4������� J�����뙩)Y�W�=&*e�-ԋ����A�!?o��-�x�ؗ���x�s!C�	�P${2�~`�e�J�(҅�����h���^ �|�sQJaz�R*gy���������-Ύ�LOg�U_��nllQU!>��$^�#���\��*C&���4+��
1�",�b<-�i���RZ`:mx��i[��<IV�|���2�'rn��9��z�ؕ�>E
��(ʲ�p���<zt�ՀQ��DSX��sy��(����O�*RRH(�}�3P�&��FkGaRL�$c�E:i�@Y8��z�O�l.K��-�ۜ��E�{����AJ��b���1[��e\Ul�:�O�sl�@��d}ס5M�o|,���lll���ѣG|����3d:������!�����uR�|�+����a1Ei���C����޻��7�}���3f�:ox1�6�c�(KYU��UaݾR$��6!��� q3i�̨��iqf�']�����a��n�͛���-�߻�JYU� ���w����g��q|LpN��"u&�h�
� �����h*�-ZB0β��F�����@�+�J��q.��*�J)NN�X+6pz��-�T'''(�;v�#m�E���O����2鳢Ö%zE��w���%� ���)��y����TB���%&��5A]��w��%>�]��]~n�g�L&�e�R��%i���l/L`O._|���P���"*�%Ԝ��F�<HްVe�h4¹\�H�H�@MR`KK5���� 
��r�o��\�g<8;ʾ�"�q���5�5-Bbzr�b!�Mã���[o����%������tn쾴��S.g�SʎO"�|^m��}��^�AeW�k|hP��h�$!� ��e�TE���d}}�Q�G<XMu]G#]�)��͜z��ʻ�esͱh:��
0��Jh�Qo]��nyl�5�:��>����E�{�d��?����8;;���l�m09����{�fY��L�Y.3�m{,<")I�I���g�{f�4?�����1׼��ŌbbB���H-��I��-�f��X�UY�l�� "���Q��ff-��{�w�I]׉&�U����7y]����#�ׯ�tp�.���>�p����c}��tzH��3�N\�e���C�ܹ����{�pzzLU5vGتi��`�A�H���hă�cbJ�G�x^!�Q��NC��EuX����Q���?�<
�|j@��NB�a}t���ѻ}����|�HS�	O�ƤU<1ZF3�/Q�����R���x<N�u�\I ;m��9��Ϭ�两�\������,����O���R�g�.Fp�c)�/ט>����jR)�(O�վ�h����%ދ%g�� �]خt���:o]�i�T&�d�£���v�.����'�ː����^`�Y�]Ӭ��Nd�MSqr�`Mz:f���;�(
��1{{{���S�z�xx\S5�`��+��ٙ�a��,K�����O��_��=�Ō�}���)���%BF��P��o�nS���$t�o�\)E����8�`]IU� F��A,Fl�vM����ʵ��'�le2�"g4����d42�QB���89z���}�R�p:]a�!4���\K����I�_�1���2�ߺX��?�?��:�,ĨX.�<x��g�]gT\[$w��2�֮!0�5��)[.���ײ�i�֐��4~-�������,������l���	�gS�k�Z(��kCʸ��2]�MK��v5&�8�PRJ��PR*/|�Jeh\���'d9�9͏�<���N���!�\2��9+���-uJ�k�����yCp.�]��191��X�d�\�Z;�L��%��9�Ʉ�d�JFy� ��j��I�n�8��5z��)K���6 ��������^b\��&��D�&Zǣ��me�mj��-�|li�2�I������j�|�Iܔ�~�Y����}��q&#D�!��uBЈ)˒���Ez�
()	�1_M1�0�p��^�����:�@�gU/899����_���H����P�9�k�9Ҍ�ӓc�}�!}�!W���h"����2��dNc�o���~��~E�����g.�\��nb��`��x_�l��p6)�Ȩ�J�ɜ����	�W�GH�qu��!j�`<Bg�|o��d���=2c��s�w�p���rNc+�/h�ckAA1!�;�kZ
�wTU���@���[�D�x��:~� <���a'y���$��Ln֊���u�8:�������J�RJV����L�S�s\�zm������'(m8=�rt|B�8�T\��E�L�g��2�� �Hcc�Z��I�=�Y�j���*�R"e!6RHʀ+�@�΅:��%��zj�Ş��;::{{{ ���T	�*��2� B�	`�~�i�7�c8̑��r5c6=C�W�itk-�'5
�R�}U6���a����畗^�,K�?}p{-q��i�t�۬�I�M�ԙ�ni�;s/:}��]��8����1]V��j�M:�"2*NϷ������$��R
緛5:G����OB�O�������N�O�=���c ����ϑD�b>�SU�)��i�b���LF���|�;o��oP�%���ܽ{����/eN�S����#v&;g�������G(�2����lN�in\����1�q�n������'6�9�_:���L�����8�D�J� �)ڌ�a���8� Z(23`r�͛7�Z3�B0�s�sh�s�{��x��!�������x0����hA�I�$!Hf=߈��Ĺ��ŝ��S��~�ƹN~l#���]]� a~7JJ}�Skm
$~��}~]���hKʉb00�毢(BqrrB�0f�d�f�u#���!�̉A`��65B2��,M���R���qȤ���h!�*�#evp�ɫ�<���yjP��ʻeB;'c��e,Px6Da��%�w�P��L�}�&ZJ�U�'�%:�R�I<���Q�3�_2���]�>�`4住�嬪�=|-��6)cb]D�ClB�'��rI=O�����
���T����đ����k�pEA��5�sG��F�v$��ш���ш�j{>�Q��Ӻ�h�}� T��ު�X*�x����g,�(4Ҥc�
z]�k���ڲ��l��?�l�IEuQ!Q�(-p? 8�My8;c�sA=A@f4�ȢT�N����⫯����{&�n�w��#n���g:;ag8�����OFL�ƃ\K�.�$�!2���|z��l���c�,c|x�Ji�޹˭[���ڿƠ	T�$zEt��j�z����mÑ��T����!��L�a!*�9D��	/(�%�@
lA\�`�O,��rF��x�9?�1�FL&4�������r� %���&3C���hF<c�L‸X1/�I���,�r�w�s>K�hw���H2r)p�$���# �V��H,�� �D�$b@����}ָ�3�!S��@��Q;Bw��5���0���|�n{�!���$�bIPK�h�*�W�*g�<#�y1g:}H�^چ|�SN�����BtT���e�(��b�S[O�
e
�R�& �%�Q!��3Bt�:˩}���=_��tӃ�(���dY����D$���HU6��n�7&j!ڦ��$8�ɵ�6KBY1���<�ލ��[����-�Yt6 �o��&�I����q�h������ ���"�k����f3vw��9��)�$(R@���]`��3�ZQ�"8�$Ǧ�J�DV�Sޛ�L&��^F�U������ů�����6j<��퉝>S��j�@	UAH��&��QV8��*z�7 �l�	y!"o��C���minUUF#ƣ=�v��ptt��cM/��nӤj���\&� �H��������~��G����˲�����k;��.��W1������$v�4������Ͼ����7r|�z!������CU�h�g��Wi�o����ۿ`>�!�g0�����,�GX.��eI�u����h{��t<��5�����y���W�\9`�J?�֯�K�])������֦_L�9Q��4�"]M��ԡahr�a��8W�G�4�lg�f��{���U�9���W%���e�bV/@�)vwǘ�yd�ne��@������< ��Z��)��5���p.zdLk�T�kc�U��/�kO�5y.@i��8"F$�t�<�2jv�;�U��p���b"�il�ZЙA��R�Ň���<O��>&̥1
$R�q"uR��ֳjV4!$�J-1m�'Ĉ�ms\�ԫ�S�YZ/BXBk�R���;�p1��λ���y�|�XϷ���l'�"��2\�e�/V}��ٛ�s�9��9���l��Fu{G����kmn)H�TQI�P4v���{��2��T*SR���u=�|�X��ƞ��{���ѻ�
#Dp��"�=+df�RB����E1�v��G�m�VӀ�bU���!5e�%�.K6�N9=�1�9`<9��uP�����-�K��[N?h1֦ITV˶SJ�G�G'R���1�;�q�Y�&h"���7h�Q���d��o�
ߑ(7M���ҿ~����E�b+wU��e �/��ߙ�����r	@����C��������c��1�6Y��9?}@9��*��\[/��s��"u�M����s�!0���4qgH 2�s�R͖�'D���;�sX?����孺��;��!���!�#���_� U@�
�'R��Uę��<n$�c�ݣ#~��[��V�ـ��T�"g.T��̝qڜ����n����oeZK"�y��-HŰ0H�	Uē:���⃇�2�)��C�����*b���$%�%F*D`A8I��Z�:^U!p���T��(0*���A��o-R�����c�Xy�SW{�]&�<��B"L�.Fh��<;OA/��L4(�Ur�$'ELNgHN>���1�!��svww���[+]����0�۶%�W��3���4'�1���>��#�=���N�&q^J�W�\a>�o�/Z�p�{�/�n���: ��ɘ�k!�1D���պ�
̞`�>�/�=Y���M���>�D�;D����2u�n�)SYJ�&L7n����:�"DWR������J.g�3�=<b��u����Өk׸����f���n�2��D*R���.�B\�~m�bv�q�C"�l�1�7�C��2Y�l��Ď3*�G:GNF�e��+�/2���:c}��kj1Fc� F���>��s��l�[)�@lȆH]-)�!�������=�����L�����{Ì�ܠ��0��鮵�婔!"�\s�3"��ݻ�99:�D�o<��ݖ�$�V]�b�h��k��󰋍6�c�����XD�P9�,�RhS�3�E�+3z�`0�Xc��ݵ|��?e�w�����7<<=&�$��S�{9���fF�*qN2f�������4n;\�w�,Ө,G��sM���yQ���GȈ1)�Y�{�Uĕ�L*���E�"ϱNPVZ�LF�lE]O1�K�RI�\L�EA`����
�R8�q.2�r������n�geK\��ZVh�8�z����gܼz����h�T�� ��#�B��1zD���3�߿���C�޽�r�Ļ�]����k���w�L�h�c4�`�?���>����E"��ߵ��گ�\����;���;==�z���A����
��ړ:��F���� |BHC@��b�O9|�ڗԞ��;�ʙp��Ѝ��P"8?�2�w>F�4V�V˖\�я�pg��S�?@*[ "!RElH���p�������egw��xD8:��kB' :�#�Τ���z���э�bf�_n��>�OLj�2e:޸@rchg^��2��B7�;������4Z��t^��\!e���n��2��{�H��Oc����6*+��	�Z�-8���9<<\ӽ�"�h!�D"AK�̥E�ͺ���+MUr�{����!?�J���{RiI��*k����R��������(�!�UJ!�GI�w���`2��4(��%"8p�ipq��5Ŏ 7�|�
_�����GGxp���3]���?����P�cM�H��=�    IDAT���n�xE�Tq�o���ɇ�̻�-�Œ�p̍Wy饗�FL&��4W�V�")Y����C~��=��KY@�^�C �A#<s�Y���H5���6����bIm�i͔R��L��2a���|��_z�o|�ufƭ�>��_���B�(W������[���;��<����
�Uհ�b�m]�3��Ղ���srr�·=����C����5��m!�5�2�w0���N�[�_�H��wN�Ex��&\�)�J��ck,nd>����I�N��.�~�����w|!v�����	t�&:tBB�T�A�����}j{bL��	�BB�2	SB�]#��!Ɣzvn��]��!�=e'�.Z��$�R�0��Y��g=<e��&�`��h̕+W�}�>ժ���,Z�.�D��k�U:�ۍ��e��Ob]���m�#l�`�d�Z����u����T�.�-��w�w?��]�:%�v������וտ��9��Z�X/��k�s�fZ����~5u�VU�b���Wc14H��_t���!il�Ķ�Je%dj`�W�~�:M���w�t:%��r�D�D��[R�.�'�6I��TyW���D@(�(�D��A�;��˯��3�p��!7���rq� W��8?=����4u��+�1�����������sL���e��Q���[�r�`�Y�)_���>�xƭ�������M�1�eXBT!q>�\U�u�x<��7�ÿz����⋘�%ϳ͜��� ����|�o�zĭwn��G�����`4d�J�@��������J/8:����ý{�x��!�yb[�PR&�h�B�и �������o�g��n�,���)�����#������_{�[��_A�@��� �4HA��פ��5:ӌT��9�{W0ِ��-Q
N>�ڲmj��`	�!Q\TU�^_�u�v�����ԕ�ښo}�oB�]��l=�W�9�R�u����-�-��sP�ր֤L�חL�U@MgS���2�H��1z���O1t�ڗ؞��[,�x�J�[�d�B���E7�ʄ��.�'b��%��s0���	���$i�Ve����墂��b4���g��}��%�ѐHj��Z���i#X�kZMδ�zo[I��2��i��Mꮬ�N������m�GR���jM �9|��u?myW���c���x���,��z���1�����S��;�Lf���z���1Bi�ƒy����P��%X�6��hLQ(!	�b���Eƈ��$(J��:�s�������k�ٌ��QK����r����߈����Fӧ��z�I�� ���_��^c�`���r5%�$":�w��SN�ψ.�O�|��-��w8<�x������7i���${�=�����0��x���woS�#E�ɖ�����<��g1e�����7���7��������?�:�u2"�@L�m!�i�L6��3Wy��7y��78ؿ��ܾ�6 *R6�*�����+<��WPz���Y��o�M���3�F��V
��6D!�A u�x�
Wo�ȵg_�@����F#��(oȲ���.��(r_���HzM����AʰY穛����:��/�3�"x�ώ�!bׄ���s�O��W�Xc��*��u��sY�o��]pĺ�#�D�}~w���n��7:���,�(����6@�؎A@(ك�D�w"����E�#j|X���a���G�S�C�'��9��P!(1�{�BJ����#{��׷6��ðvH:G��,"H�ሽ�k#\ erbh(˄1��6��nk�\v���LW��ȑ�#�-5u�nFD��EI��庝e���e�ēX�p�6jO���ڈsv��KY�����A8}�sk�{��*�n�O1�I�g8פF�Lᚤk}��+B ����x�͂I��A`2��/8�M�5�
��(�:�mf����HH:�&�_��8�5f6l��TЄvSsM$7��!���䭂�PJs��*�kN�Θ�N�Ww�yx�Ã�P�h����jQ��FF�_�kO#�EI��:{�Ƀ/��c��9�����������?��]��������8�B��H�(����X�\A��������A���w?��)v)kO�z8$O�"wv��wߢiQUMҝ���f�NNg
Q���� /2��9Z)�,#xP�h8�ȇX/�JB�$U.�w<�l1�G�lW ��mCŀA> x�=8�瞧\Έ��*�*P6�c���e�J%]�G��5���y�����.VQ��6�0m�O�܇�tkS��^�\(����1Ɣi������3�jB�!��R3��-R̤���<���?�?��O���+�R���e���4������j�r�RZ'-�NU�&�~��&V@ˎ=U�\���v�%A$��PIZ�5�����&+��; �8���2M��ʵN�G��n5{/k��;�}��s��Ɋ�H����}j"I�ä�a�j��!��/�[���b�.Cv1&N�~)�"�;�����6e\�"����Ν;��x��g���4���3�s���>�T.�]�wL����>���������>$)ѕN<B��nQ$�b������Ae)�!Yw�^�ʲ��:3�ImBH��&�� ��wB Ed^V�,'8:;�t6�iB$���b��p���$�k�Z��{O��Ɣ����-o}VB�;ɻ��I�`�eX<&����ٔ�����6��}Ϋ�(�d����>É9 3a�г{�%n޼��sh��46�E�x��`1���ѝ{���_��1]���`=VW�y��}�`�[/+��z~������-��9�7<����o�����v
$�dgr����)�,/�^0_�P&������cr��U�`r������hYq6]@��@�Vx-��N�.Ғ�w��y>����旿�%y������b�Kդl���.�:���k7��9�iq�����x�`�Z2��������֞w���_�;���]VuEVYFӤ�%�b<�p��Unܸ�����կ���Ͻ�p�qxe�����V3�R8�BT.dĻ�;��:5~�!]�֮)�֙�6��>im�@�{ t�C���u��.��e�������>Qs�9�:\��{C?�fah��HL�*�t,]0�g�iD�"6um
�����j�T0��� O��?{"��j]�s9Ep>z��QH��A����8��(�E�ڢh�l�ƝgKf�����}�$ӻL&�����,�+�!�QjHJ�z۪2�-�s�Zo��.ӷ���8]SDb��Қ̨��iA�En1b��`P�)q�rBQ�F��d���j�X�i_҆u��7�R&���p�^��uv/e(?^r��e}m���؏����?����M��M]˛n�� ���qHi���̴�w*�����[7�w#D�m`�/u�$���rU����w��9�fMC����v�I)%Zl�Mg���i��������CJI�$AIVJb��2���i�����F`C�ɑ\�Nvp%ӳ�Um��$b�sD�L����Ղ(���,�*GsAm��d�g��R����?{�-��ʟ��C����O�ۿ�[>8���4IUF	B��w�ի׹�ʳ���<{�r1D�{�7�{��^x��_���&F�C��@��!#�)��y�y�կs���64��,8��dʉ�(����'/,1��u(��)��[������W����LN������D;2�Ny���w��ZK����x�eȇ#�!"����g'�������q{m�,ؿ��}E����Y��,�J
��w]�����C$:����������b n�5�������i��-���C�R�*�-�K����#�'o�^�h*�(D\;-���!D���@�x9��B����_�1�D$�@���℻YN���s|������������x�x��;M]R�UXwe���EX�Iڟ��c]��=ן�J)��J
�4dENn2|41R55��$J H����qC�9}��uqx�����9��x�~�:�Ɉ,�Ę�SG�/m\� �>��!��E�>ٹwc��ߕ����9��f��
��0�nC�%�<C�5���q�u�y��y����"����J����j[�^g�c��GR�����Š���\F��T���L�04,WV����5���3�v���!r�`MRJ������Tu@G�S(C��b`~��;��z��.y� �5|>�˧����\�k��&�n<��|ͽ{�����G�߿�(˚�jh|R�@hL> ��q����u���%7���}��p���ܸ�?{� ���{���)�]�j��g^���9w���W���4h-[8�!D��Q&.��(��Ӗ?/�_^V����_��=|�6�|�@��B�3CD��<�V��lJD'꫱���L��A��~�<��V��.�-�'��n�e�,x��]t�.�/��J�����k������[��o�ɤDH%���k��я~�T��Ȟ�髚+"��EAĐ��ZA
�]Kbk�[��µD���'k!"	�sOF���h��s�j�o�x�����s��Y,KWS�U�4U"�\��&�`��,C)�`4m��M�[4�z�i�n$}�ņ�9l]3�(�K�LF#�Z,�d4�v�ȱ�>6M�&�����E�q���9����}�\��0� �+������r�.R�\�*u�_��u���c}'���k+w���%�&�� S��V���µgO\g
A���L��A���(|�px_�뚥�(�ϧ��۬�vA`g����}(A�w�g��甍�llt��Ѐ4�)(��;=!,O8��M�h�9���wyNe�H���+�-.�Qx�8Z�yx^��Ś,����p����C��`�f�l��L��QJ�1%	���J~����7��_3;?&�
�cq�������d~6���y����׾J�<����89:N�6F|��4D�� ���T�^|�?���y��w��f8QV�$�%E9-�xޖ��ylD�{D��Q��*lY��d4��j���$H�9R�hr��8�s�΂I�S��9������H��ҙ����i������]�8v��u�����u��e𕋙�K_�A�bh)�D� �U��Z
IPR
���R*ɤЯya��˿��ŏ��/7U�S���)2}AHQ�c�QDA�!D�Iʑkl���^k�u�.()pw�12E5K���)����W���=�����n�\`/EaA`L�p(�~�()l:e/frB�(�����s(18��&�w!A&�#%"�V��i��(@K��
-����[,TU�sn-�V׏�jO�uYî��{鵍��Ŏ��ǡ����vI�r����u��~8��l��A�ׄdj�%�Y�]I�����I�Q��J�nJ��9���!�+V��Ya�%מ���4͚���%�si@�yY?{��w��(|ʸD��5e�����^�
����3:[�%�����ūe
\+�pT�(}��5�l�K4�[�0�K�ǣ��h7�S&��^�M6��	��g��������;w�cw�">�4M���Q�&7�����;_Q���������q<����z#Ā

�2DTT�����,=�p��n0��?��?}����6�H#��k�TD�Jj1�ֱ􉛲�4��M]!�G�$/3F��B������f�'b�� IXJMҠ��B>���|k�ɞcwO�џ<Hl;�k-��!`]�K���8:�ʶ�ww��n�����\Ƙ�|b���wY�.����(��h�
�C����S��̞h�ԶNٽ�VQ pi�ƶ'���=w�9^��:\����������[bg)�"��>~x��x�`�q��3�	��ٛש��:[2�mCpĹM'U�	�w��~�i�JY�N��{]7QzD��:ӧ�a4`�%�e4��,	��(������lFh9�V�!F�њ�>���:���bЋ�z@�$�-��n�J�� ���i}��Q�sS����uI><Ew�!D��0��q5Fzr�6�P/��S��/"MU�Ɗ�1�>��V����od-^ꕧZ.��\�ju��ޢ��6�,�kb�����TW�o,%O�e���d����>68۰�M�e�29>"d�!�Т9<G�S��y�:�gXh�sc4�h7Y��������]>��`A��DR5�5��p��-�L �%Kp��^$�d���AX0;u����
�
��b��IE�"������� ͐ݽ]�S��3&;{|������]�y��N%T��T
h$G&'�L�J�J	�J�F�Nv\�W-�MIaB8P�Lf������9�k���C�ȇ,�%��]�Ԟǁ��NT�v��>V����`�7Y��z��3��ه]t�c�;�n]�	��˪�� �����-���)cZ먢���XU�(%kQ6'O:n�ڗ۞8� ��1FA$��)7'.����.?�%Ȕ�=�{�=Q�I�	1�K��6C(����ŭ�����7��7��1���ӣ����`�)Z���
����t�����u�|� ppp��k�о��r�!�ј���6�u�b6Gg�"��;�gw��Yܻ���(�+>:�s��ݵ�v��ԕ�����l�'�.K�}�sc����MRlH@?/뎫���/�eY~,��]VnY�V�.���w�^bDӠ�F��5��d@�2�����`?�1�����Y�is�H&�d³
5"�(,Z��=�b�=���qk�ZC�L����������ن�G�޲'��{�#±ZN�)��J&٘���E	�Ai�򎲶(Q0P���t��Zy���<{�G�;?y�����ǈ��/:�oU-��U���܀�+f�#�� �BD� n��,�MI�a�*,��*�d#��l*�
0BcИ�V+8*ϸs�.Y�QN ��s���}�޹�u E$3���[�wIV�%��.���k�R�&`P"�D�u�k��',�g)��=��2�C�6�(�H�R�,Ǟ{��(i��~l#G?��R��ہn��w�)]0��襱����w�)���|�� :�����]2�;�~��e�_ �n� :8q��&�gY"�њLD��VRZP�������~����O5��ڗʞ��T �S!2��ǰp]��9"@�D�Dۇl1S��6JK�.Q���j������*��_��W�
��3N����}����M�HZ��v��|�����Xmuõk�x���y�7�˓F��������c��%�n����#Ƥ��̍���_��Պ��������5�=�u]�컒rw�Qv<r�.d�>.��4��uY��(1���,�,��yX��e$��!��<Ϲ��Vg��9?Ƅ���1��Q�\;U[�shR���cd``!B�ȭ`��ߪT�Z��uR�h���!��A
��
-FC�IFÌ<�,����Yׁ:�[�����w-�sY?�ݧ�cAGr#�(�@+�tA)�'��I��̀I6b'+0Ab��AU	4o��!�E��C�%=7n� V�z��v�l�ݻ����v�"��[����/؝I� ��[[�����,D��� :3� ��(��ِ���ͦ�|!<�Gx��c+�O��g�����W_������������Z˝���|��I��u�ٽ��#�_A�֝�B�~���`$����2Fv&c|ԞԨ�<QD�V(�m�4!9��e��)v�'[��ܔw�������=w���q�6�J�-��u]?R����9u}E���("��>����Һ�r�J�bBD�1AX���ڷ~��|�G�	p��/|j_z�T��Jʳ��� �XDi�@o1(��l���2s1�25��o��h�n�pas��	�T�W�����~x��O��w��htH����]BsnJ��|�(��e�p�A��FG�"h�Ŝ�#j&X7��,����������c:9Z���j��ko�91X~�_���Q��|t��[�'�L�.{{���M>8�aS�L��`4(�Rt-k}�6_�R=z7���"��Is�����F��E�923    IDAT��a��}"S�3NΎp��DIUUH��T��\\t����b�ɠo��1k�f�b�YӬH)ט�>���]2� 	a�d�TPާ\����.;���+��L��>��3�R���f8,��&��K�JA-�2eHQ!U3 �į�d��k��פ.�4JR���Q��s��m���Q�^��Mb]pr�a�ƴ9c<�"c6?E��h4$<��8˚$#dMN&Z
��1��2)22�/���+��2�p���W��F��#��+��E݀@�0Z`�@���9�7w�B[�젅&�	�J�5-�Z"�Lu�~�Q�aA,-f�!W%�mL0����Ƃ*dM���iSsH����
�q���˺ϡ?�y��g������\Sw8�{��BF<BEv�y�+�\}v�`��w�l8b��ϲZrzr��{���w�ِ�%.�Zi�p�q���K��[����|t���������o~��vd�{��݆7n������Fh2�ϩ��9��x���P7'K��x������9 y�*L�b�W��jB�qYC�A,MI:qa���nQ��<UX|c�9�҄�D:�S��Aw�� X*��i!u]SU�:��֮��4Y!��1M�\hvی�D�w�k��U�v��#�������{}|_�XҳWkk-VX\+'���`�@{7'���$�r�L]=X�b0j��"E�Rx?�<��;����})�ɜ���2
DPA!�"&K
�պ��I,M� a�l�Ǘ��t~�B�X�ns������ZK�+T���d���]��%?��O0&��H�mp�rx��׾�7o^���!���|�������p��}����p�����l�6����stt�l�@J�.�Y���Ų�xmkC��z*�oG��Z��9���� �m�*�׻W�������E�:����-�~\y�m�AĔ5�ϧ����;>>��ÇX[���CYm03�g�����MfX�6��:|��V�*8B��hR��#ovM{��3'M�0���4y��ޟ��'L�Ӥmy� 	��᧿��B|�o-���1�=��2�����߈�����l;j#��<u��m�j���V�M��\[+�9E�>X琤�R�ܤ쉫+NOO�N���9�o�f>�o���,ţ|r_��`A& ����K���>���|�{�s��}��!U�� �@J����(P�	USR-�9;�����?��)�ߝn��ҟZW-rcȔ��Vܽ��Wy����وJ|��ort���`h��Z�)��1�N��he�-���˔�`������6ӿ[�- j�EB�J$JI�4D�xj���u��Z��mw㷿gte��-�\7�
�1$R��֦.�|���ϊ&�Ͷ3دh [N��t������0��	�bww�3V�eY󕯼��h,��yQ�Ri%�R���Nc=-���g�J�� Hݺ1����7��:�3�ݜ�v�g�  @)����i�dQ����Op��k�(<�/O��j�*�%�-�	$��>3��v��M�9�ވL 3� $쵀����i��������	����y?g-�p��#� M�`����F\I)���?�W�ݼ�c�蓎C����k+TU�{����ﰿ����s��9L}�� ����X�vv�������]�R�����C~��1<�X��˗Y]]mnސ�a�댛뺤(�MA����O.�>���	�/���S�p�9DS��pOR�}�c�puͤ��Z#��p���}PN/x��H����pt�ϣ��2���.����)i#�ik��*�ڢ�	B������nۻ�plx 
BZ�����5�W�:���h�r�lRQ��Cʲ����0����XWRW%Q��R�ѓ���<��K���O�8sp�ǃ���#u���6��IW�����Z]Bb]՝A������r���p#�p8D�U�4F��\< )Rx�18Sa���y��+�(�y���n�b>�#��T����.
?��צ��>d,Ǫm��£�D	��,���z������7^CĖ�9i�Y��*/*am�kCʣC޻�BL�B"�"J�$��V�ID?��#AY��{�%�b����q��W��M��O��n�٣�=J;"�P�#|P�.S�_��{���7��N4�*���I��c&�!*2�P��l-�鏮�]�+�څR�m�.|m���Сut���Ű�!�|A�9!�ɹӴ��/�n�Y�X,j[��ח���p���������`0�,k���)˒�����W�Z�����qB�}?��sc�'���O�������b�}9>����H�,f��%�ً�l����Xw[�H��^�BI8�� x��$	:ߐ	�#�5Rx����R�q���W^���+X[����-Y/�Ҷ<dooo׮��/�@��x��{{{L��N��-�89�t�C���5���Y���0n�m4�l�2���i��k'���,��l��$nM����i��^t�ߓ�	��{��ߦ�O9<�G)	ޒ�9�p̷~ɀ�!Hw���4�}C����Ǐ��ˊn�,�l<�p�5oj��`m�1%��Ԧ`:�������!��״���ԅk
��)�?a�M�ע}��������.yp����Ģ���7o������9���������
�Ǜ�� ,9:�FɈ^?�dIg��Dw�4��x��MP���Bx���.���oY]]����<xp?,^$S7�U���00�3¡U�	�]����h����Wōb�b|������|F9έd��t���s��w��}҉T1�%�T�\������B�����&/�>ZG��=�:bg�����l���y��"�s��%Dg�&>3�z�5�u5�G���Ѓ��Ak���ۚ<ː��L�@i��e{����Z'��_�)�_+<k�4M�� l�R!�h���0�
����d;cʲX\
-e����~Y��n��k����&�	���
����g�g��ё�L����F^:Q�z\:�+k�a�#�/�w���r�,�� ٠e���p�AVJ��ټ<e�Z��l4�[�;�B�׸z*�H�H��ш(�(˜$������������C66W���g���3�������e>�G�[��(��#����l�SI�0)k�t:�$�D�0[�Z[�ő\>:�ǡ��^J)ZT�S��|��Ok,�
=��]ݿ5B ![�k�̡4�������H�g�)2���Y_��=��pM"�r��^Gm�(B�A��£A�T�u֕8_amIY�p�0�g���P�9u-:�x��΢��8��찰[ �$/N�s�=<s5ݢ��t�Iӌ�h�$I������&:D#�GuH�1�4�H��a��h@��U[$Ƒj����>��t|�/���q�����	Y/���R�z)e�?��|�Z�
P1�&SY8��Ԥq��2�m�����X];ǅ�A���%���C2�IJ9?"�,YoH:ai�JŊ(�w�҂~��f�Dc*��7����(���7�@�����=��#���^��hfӊ�k{-�"���h%I҈HKr���(x�?	uW�H�k �"�_0l���4�n����Py!:ZBK%i3����5ݳc��l]Ҭ��)�<�\#fA�|l/�
���d7oE����@�mO2��������I�1�����a0��?�w���?�7�@J%�?U�����+�|GR�U�g�z�ϻ�����~r8焋��	�����^;V�=k�\�=����c1[.����v/�i�l
*�5����`D)f����cl�o��7��u�y�wl?z��!zK�0���!:R	���p|r�`�#Mz��c�8���Q�5EQ���z=&�IW��� Z�(Uw��{�@/�!�F<��(�$a}}���-z��P/�(._;�󷼂]F'Ϣ{�{�%;ۀ���t�a��q΄V��x	R;�ڰT�6+��O�kF�DhW.���]��7�� �X�\�?	�(_S�I<�U ��B8�j ʡ��69y1k��,���Y�5�O\��2H�(�)Yo�J"�bwߦv%��,�(jKE\�x�^x���M�$��
��ίG���H�\�t�˄βGH��)�����"��;��5E9eZ�C[Ζ� HQU�z>-B��#�'���k;6�'�
t�$��XW�d�d|�/~�S=�a��%ta�E�#._����\�r/"� �f��;h����R�,�x���'K&�}n�>J�X�or���Aµ�����(&������dDD$:
h��p���\Acp��eLxk�!�z��by��z�E�vQ�=+�m�s���R\�����ͭ�W�u�֓$a���Ÿ)�H�p��.z��M{��\ӑpg�ݟ�tY�sJ);���xZ)�9:<A*����ß�ٿ���&k�k8�y����|�����y.�2�x\���NƫZ��*��y/�/�{<�cC�$�H�{�Cs������ܾw�\�]}T;����27�)���KE����4���b��d��T3F�>[�׈#���ڵ+�e���;�*��K�$I@h��G'Gd��,���$I�|̙#�t�܎%��
MܗpMK���-��$���b�z=��{KQ��,�����E���#}X[���^z��Wd�\5��%΅8*c�MF����~��qO/<��+A����f�ǟ�N!��E�bm��AZ����Y%]�^`�����Bx��g,x���Z���эi�j�oQ!@i�w5:��y>�xC��A`a<�~�˗�r��u��~��*��)��y��:!�����9�PQD�#Ԓ�H)�ܕM��7|)C0��iLU��"CHRTd��ȃMt�/,Z��s��N����炝H/I�.��zNGr��o�����h��G�$��`��/��*?����À&'}t���T�Li��V�R�,���S	�e6�p��ۤ����&�%��fl��1�%L��G������;4�}S<c �|>�4��`d�MXT�3���`��8��>��ܙ4����	�'�
��3�罳�-����P����8f���M]��g���B�ݽp:�m�����p����$�e����U�慗^������޿����E����l����'T�%k�ON���f�p��o���ّ���������8�� ���|B|\����y��&�m��l�p
-�
0��:�o':J��)5ei��=�ш^���ã=�6���~HQ�Y]q|b�N�E�x|�(.�
{>�vm���SJ��=��RW�i1ĝ�_�<�b1�ڬ-�<�ǎA�HR,��Hwj�e��PB�z^���/�����f���l�c���
(h�w�E��ؐ�!�,P+�v#�@���x� �g�>�pq�R�A�~4�_���_��x����	��U���(=B��Ƙ
c+�(%I�"�����-U��-G�$�X<��^�|6�Z�"M��DQ��|�#U�4MYYY�r�[^T���yM��*�D��'ME	TEG�B@)��u�#��7� )ΦAJ�Ғ���Ee1u]1�N��dYFU5|�S��pm�?�L��o�z�	��H�{=I#tB:��b�!N��g)�����c�jfv(���o�k��X[���
��#Bb�R�q!=RA�UH7�X�� ),G����M�^����*����Wz��x�T�y�uQhѱ<ϙN��u�Vqb�Ž�H��w���{\�pCגn��)��Ej
��s�2��}m0X�\b�����9��.E�U�.[��������i��M�|ip�m�T�<���SǱJ��������o��K/����XҊ���ƍ�z=����r�
����]�u]+))CI���[�[o��%��/d<W�W�W"�8a�qRD�*�,�cP���^�����G�u]s��e��~C`?�����4M?���J��O���2qj=#QAҴ�wtF
�����]h��Q�h4"N4U9�~�cv�k�����~IQ�qƲ��M�Fx'������3��9���\<�۷owh��񄕕������_kݥ3�E_Pg��7��9ٴ��ޓei�bmN�)t-;��0!'���!�x����*&�6���>��g.�s�>lϣo#�AW�5)*єEN&EG�|��V��!��w U��-�=���H���a4�ĺ�JP�K����>\���eN�X[gZ�@QU5UU�kT,�O�j���>�R�����.r"E����Ue���e�
��������}�����+_y9�9ͥ����
��/��n�]��BX`���c��L���2����3T��~kmC���������X�<���a�W�K�ʃWbʺ�zE������c�X��:!JRfSà��&�	i��%	��q8�^�kV��^3�`��]+e���eN:L��qrN/Yc��}���?!����_�7ڢ�'�B1�b��.8hqc
�kx�H9VVW�(�g�4^�?R�4ee�����:�'3��)�+����g�Bт�!�[�����,K⸇֊�*O)w�E�֚���Ά(̹a^L���ڊ%���`0 `41��-W��W�!�i0���NY���c�$ass�[�lnn�2ڠ,K�޽K�$lmm���#��9�� �����ϟ���<�y����w����Ue:�<����>��6�����R3��.���(k!���j\��[o�u�c�_�/��x1l��.rRJ��!��{!�Ctj�g=����p���*eYvR�4�U��SѐjC=�lo��@D][��7d}}��QG���G��,u]��:
�#��xb��H�&��7����t��YAQZ���7���[ᵫ̎ /%R��Izy���B���e�}k�ܒ����/�h;v�N�[~�?No'�4MI���F9�������v�פ���@h�FQ�Pck�
��BL)�����q���C���gg��'���/֗9o��k�����V.��p|<���)%�Y�|>'�Ť:�,g�\�φ�c��*7�%*��%���.�э��sM1�	|�Ó�o��,��g8Ҵ�Z�"beu��h��|ʠ��7G���(퉵���3�X����h-�g'���?��0�!R��Sa=�C$<�/r��98xȍ7�<_ya�A�`�D��Q��	��#/
��#/B������67���!/K�
��F*�$UQT��{�a4X�_��&�^�m���t����;�YƬ�hP��e��cNM+��L����;w�<\����j�vk���v�P*�R������0Y���z�M��������
��x̵k�XYY����{��Q_�����׿NY�ܽ�����,���{ܾ}��lֵ��c�w�9��\8�R�ⱃ���g=>��#����(�9'�t���>�Z�\~��ڶ��<���ڂ�I\��c�p=��cyH/�v`}/jՎ�l�����q��9VW *lUr��<�WPy@��-�4%�"VWG� s6�6��v����z����!�������X�"��-a�Cv\k	�ϬtR*�q��vZ�;��v��E���,ӳZ��X����+�jS+I�$D͝`�A���l��V�'��h�Pm��2V�p�!N���uЃ7�0��]-#�tqv>��}�t�d�?��%%��-m��f���6�Xou��s@���&��3��L��j�v�U��B(�X��u
![���"�T��M|��Zy�%���p&��,�B�H�n#�~�CE�աɋ�8θp�*k�[���*
����
c
L='�)�������_{�e���]��<P�Q@[#�p8R*��J�DxI"�ق�b�g>+y����%��ӿ~!�H��TL*��(ͨJͬ�QQD�E(o�r�:_{�޽q���Cjc���'%�� qD����~�+|���y��5����c�ݽ�/�s�ܹ��GO?�˭�v�߷T��(�⮋����K�\өq�u}rr�xr@�e"�)q�q��Z�|>i�C�1��x���Q������p���z�%;��Zs��9��kkkݜ����ŋy�׸t���ܥ�-k̋P�~��_%���w�yYS[h+:�Ҍ��Ka��3!�!����e������+��@��{JJ�Fz�!�    IDAT�{�kZh�����c��<�>eY�]��J�i� ���>
^bNڮ���dx#�d逵�67G�R��!�uf2p����F��3�i����e}�!i�����pttDY�$IF�$Ե�"�Zr��-Ue����C��Xۺ;�SEA�&��hbA\>Mv���RH6"�� g�zZ�x��
=����E9 �M)�w�)�C[�k�@�7ކ�)��)���v��E�v��:�v��`Q�dԠ{B@��=X���<u(���R���EԡގP.�S3 䂪�Y_�`}e��ׯ�#RM��!�7{ё�E���+�ٴ�'d(R�u�s`}�ݮ��6"�.�~���"k+*Sb�'�R�b���׿�������g�lz�|>�N�x�E���	�ϭ��g|�O@I&������ܹs'x�	���x�w
SC�N*� c+�g�d�`�;�X6��Ylr~m�ee�ޅ�T��NҌ�L�����4����.���}����<z�<�69��A���k���:���&�뛬�mP�5E1gw������?�1�*B������D��A5)0����ϝ�E�ϟ�d�t:%�SVWW��stt�TS;t$I�^��
 ��1�O(�^�h�JU$qF�FL'��N����s��9^x�&�	{{{L�S�1dY��/��w���R����|pg��/�e�yAkVVV��w�y��n9�a��B΄RR���������������/d<�zw�Z���.Fh'b�E)^
�&����1g�7�2����jUP�;���YV�N����>���.L���*[[�����)�6�p�2�M����	�X�,�ܔ
7[QT�e��G���<x��������'�s�$aee)%��PH���[�!���W�D����}ʘ:���E\���!t��8�����X�7y���BȝQ�6�^�cl~_iI�e�#}(V��(a2�
'�Kdѫ`� !��#}c�,�`�9����ؠ�E"t��-Ri��o��A�#E���g�������O<�X6ŞpOR���"HVV���7�䅫W��S�,[��pO�:�d�T����ĲD��
)u���'�"�~�l��l8�A�{����F�1��i6o���ˊ�����]�_;��)��/w���<|p����S��#��6YY���7�/}�Ud/a:=$M��}�������Q�BH��Y0zd��R�%��	�	�h����1DB�瞻w-�l�Qo����YJiJF�b��T���jDl1N�Im=�2�G+���-._�y�c�y>&���qJ6�&}��h���j
��>�����׼��;��:j���S5��Bt
�6�m���pQ��-�~���z!TJS��$I1��(Jf�)�露���{TU�����\c�CɈ��sD��L�ۖ|��Qy�wԓ6`8���	��.{��
R�e��W(���7o��H���q��^�=
!��H%Ơ��
����2���k���DJh�X0�}��]��=�}�����$鐦��i��5>i{7�nИw����H��b��367.p��UVeuL]嬯�S����f�&����Ƶ=�1��U�(q3�����`g��,���*���7��q�"[v�7�4��c�E����/��j�Ek��i(w�vN>��h��U6��SzM�P.dAl!���@��+�� �B����}ֻ��N_*B[�
"I,.\���9�R!�-w%q"�����k}#
���e��G�!�
���]?�}�g7�yE����˺�Ը\2��ڵk|�+�p��y�j�mK8��L��k�m��k��N�nz���m��YxHʈU�E�DIL�H�>�����E�aHe9�������W.l���`�5׮_a2�g:>�*J��D:c�_ޡ�����X�(�G���������h)0U��B��t:�,k�h~�d<g���$JgX#��!��~�w��Z��n�z���&�����u�ԜL��Uh#��"d
u����c�pD:ec}�nUR�S0A|��2��r2�b�GE1eY����O~�c~���SU����i��\���e��5a.˒�|��w��҂{mm�_|��xʝ;w ������A�M��$I�1O��ʾ(J�
?��666�R0��h��x����8fss�8�I8��=���tH�ݻG�\�~�<��ƍܸq��vm�]���1���766��o��eǿ��\E_m���v�:@�@�RI�r"���=�[H����8[�곎���}��]�:�eMU��<��y��@r|R3��p�,;�����\�r���5��)���[��r�w��9���ܽ����}N��R��X]]Ek���.'''$I�e����J4����*���->����=^���O>���w�����+�˿п����Z�F:�
�X(�������</B�֫���@4�7G@��V�L��;�s{f�p�$����*��ƣ�`�ӝ�%.��is�������Q# ��g48T����
_׃��3�c{{�|:Ai�|�\W�i)�.X	}�l���i�K�M^P�j!���DЅ'1^���ț�v��SCu�g���w皮m�O]��p�&/����?o�ƛ�s���m���>���Ջ\ؼB��ump6(r��)�uă!��~����o�����G��\;�xf�`:�3�嘍!�d{g��}��T��e���H��*���)^&��7޻��`�H������?���gQ�B+*�8>s��
Q�����xj�+�tD�`�lBR;�`o�����;��m���YY��e�uIU���no��`��v�B78O���H��TY�M'�/��� �K���8Nq�5�^AQ,l��:�&M-i1:+�V���y�3l�ᬵ$I�����C��@����=N�˂��u�(���9�Yjk�D�&;�3k;E��я���S�������H�sBi/�PBJi�.<8E�mbiE���K)�!b��z�4-s,�g<O{7��<�D���;�,KI{0��u�����F}�^�ʵ�3�N�˒���]8O������׿�-{G�$�ek뛬��1��893�Y[�h���[�Y���K�e�/�B[�"2/P�Ӧ��b!��=�����}�Gl=�
��m�h��"؄���{iz�$�eKhLӚ�h�q(!2�x�bmMU�H)�W��s�7�7m��\�E݈�G�%�?�aX�-��|Z���'��%tԇeN���oݺ���#�8��s��Y�^T�Y�	�7�\
%�:>p`A
�p ��&Dg)�2'�ׇ֤i�S�e�d2�,�ywjۄ�r��4�-P"�ރ�TE����M���6FԦ+��xop�RW)��u�DhE]��������.����gS�xE�:ؓEX8V���CƓ�y�P8g"�������W��[>�����VV�ܾͭ[��̦H����3�Lx�h�������T6�c#"G��CV��,��	4��䓒[�n������?�Z���j�zm�"$������{�庵ܷ�a�h��s�$a6����o�����$	�����j���eMk��q�z�eeYrtt�|>��_�Z�I�0:�s2�t����ۦ�lmmq2S�y�w:88`ww�?��?������g?����.���B:�]�p+�l��/�?���E_m�L����9Q�8V�>ʍ���F��DG�<�i�cpQ�	��e����`�P���sDh�Z'I�U���N#�	 Q*A�cBJ���j����Rtxd8�_^�M��y�wv�ȁ���d����ܻY��"�J�[�_cw�psJ��q�ҋ\�t�G0�?�dg����M67C+���ܻw#������k��1�s|r���Z��"�S�ӥ��S��Y�m�kreCFr�1P�_���&Uh[C�C��d�MVd��|H}BӋe��Z1O+��OA� C&��|�><yq��ƺ���I< R�T�GD�,`j��b�^�#6�]ccm�)��cU��4R%���c�$l�X!B¡���%�[ba�eN9�G�>��H�^<'�%B���S(J!�¢�EKA�<G'cD�%C&�l0D�����-�Z��Y�׶ЯT�����H�P��v�pB`e�P���H!Hc�)r�|LgX;d|,�	����9��l���A����`��B� pr"B�^���+����r�zN;FIƴ8��H�r�2#B \N,���)uY���^�э�Z���M��'�~�uQz���s�QMP�` $��}~��cNv��Ͼ�o~����$!���%Η8�k�7�y������_���Q��}�V�z�kN�czf��dʃ_�7���g?��ܕ�B��З�K�Jcs�4�H� I2�x�w���=���>'''�'B@�G_D������� �qK7�AtH���:�^Hp1r�����#}�-��`��&ZW7�8,��eG�,I�P� ���ׂ���4�ac�!<��
Q�'Ix%��$�Mf�	u=��_AG�a6-H� ��)�+�p
8B��`�'�F+8�u����35�Tp�Σ�$f6�09�Q"���P�N&��"�bp���\8w��sx`0u J��yI�qIQ3!R#�Y�)2� E��;?N�'�5����_���я~�I�޿_���E_��;m�y!�x�W�[��y��Y��
�۟����a}-��JRX�����w��������"J��C�:��k�X0�������Ehlmm�ꫯrt����i�t:����loo3���hD�$lll0��L&݃��W��z���e,�-O0�?�W��/H{����AkL0�n=c���X��$���U.]�ĵ+�Q*ؑ@���������{�j⤼k�=��FKh�0u@�A%8')�c<eY!�"K��C����A7f-�8d��U�)���p��s�a��G�P ��� u
T"I����Hc� �h�k(~]��@zZO@���X,"�'�8L���ru�{�N��ZŌ�#և#�sN�w(�YE�k󳞌�2�rHx�Rz�j��;7����o8�"Q�%���5Ζ�C*�������������%����Uf�O��O�͛�(����n_�����K�c�R�RAY8�u�S圌UY�_��� ?���
\�5v�D�T�M��+���Ռ�*��>)^��-Fh�6�[�:�D* �
�-��V�I�`�
g�BL�1E9�*U]�l�=)4Λ`g�O;�V��F���c�ܹ�p8ll^���
NNN8::��իH	q��c�ֲ�xo�L���P�U������Z�S����0���oZ�WF�QE�M��':�_�/�x��#��JL�ｗކ�+*��v�mզOg�C�k�i]z�rw�Σ�Y*�"�x|���3���ˬ��o\��>��`u��x��ct�cw����;��Q�
V���[k+\�|���-�s������n��޶��� ��a5ݴ!����=�W�l�v�ǭU���j	���������b#L�j����A4-��[H8O��|d����ۺ���E9���T�	�m�k
i��Y[nՋ�M��R�(�J!��?0���d���>��P�B���I��R�$��X�	�����I�/]��ڧ޼gc�����6�]�h���A4���*1¢��a�����@^�������2�8��
��"��rw�*X4"��� \�
!BKLـ�{B��V!��Mr����{���/��M�^��)����ȝ�ߡ͚������O�̇+��"dDGo���|p��7�)BJ�g���]���������h�XOY�sgkL-�#�3��wnq�w�Z�e}�S���J$D�	�����{�K�8�RD*9��Ԧ��΃@u����A�-=�m�89��!�2�V��'�^�w��8��K��ҋ(5U�1�ƒ	kPJ൦��࣮J�8B)��hN][��5��'��TU�3��P��JE�klm�u�q5���AG�Z��f2ws����$x���EenQ2�ʕ+!�c���l�e��r>X"9�!�C)���D����U�EZ{]
YW��*�s���e�VE���3��\��{v���HN�"M���������o8?�����V�׸�R
Q�������.��qtt�W(-��bv�<���f3����`����k�G�8�"��޽��Qh�dY����Y�[O"з����;����4?��?a�Ҏ�3RH)�|������;���>B�< �q�R�5'�)�*q�P�-n�D	2��Ea��z��������=�$j+�k�����}*k�+�s0诒d}��*np��j7$SHLT�E�fߟr���=,l~�X2�>���$�)�Z���DR!��U5UQa�G�4��p��iS�36l�w8b�p�" *a��8A"p$�uH,J���օbNhjkR��y�7���]���g�c��e:>��WDk��Z�|N�,C�Z�6�u�,�����!&��:��U𜌢Z�]�0t�`"��KZ�4E�R��Q�,�b�>j��Z��mv���Jΰ��ƹ(�J)��!�E��`	~�����2�rh���P�8��0��\й,<�8�i�"�u��WW��RjSrr�d@7��$�J"EP𛺤ȃ�6�����c����4~�g=:RX[c]��H5�3�XF8�I�OӔ��5z���T���u�]�v�S��(�Nk�ׯ_g8\��������ˠ_�sNHD^?r�?���s��]�_�/��X1lxo����ށw8����[ŧ���0�^����mW�4��n����$Iё�*s�}��e��䐣������>�"1V����!��`����d�ݻ����X���#N���'�F�΋��r�����{97��� �g�E���S/4K�x�����޷��l|��llm���m6�%�f��W�d2~�Vo]�����1��cY�eY6�����lk�[/qޅD����N�m^�0�����9�{�N(+H��N1UAU���\Y?���*[�xW1�3�}�No,^�<�gi�x����Q9��:���$�ܮ]�ֹu^z�%F�!�*�{���7?@��Jǚ4ӤYL�hL�֠T[ny�M�ƅ��&� pE��;�u��!����|�B�Ƃ�2���X#�2���Ο?O����p�i�R=��S���G�C[�Ra���!�$R1+�Оs�x���\ݕ���uU��yn�nh���K���y������siKyP�1�k$�������Q,��L`G�"�r�k?$�!d#l*�X��R;��}�rY`���8g�Lf8<Q��T���4�#޷Tp�P�s�*u�J~��!�Bk�X1�0Gp��a��$q���.%G���tʅ�h�%�akѴ�ei���̦ަln��_&�2���!�E/�{����[�ȸ:��ϻZ���i��U�E�H�z|����g5�nˈXˇ;��O�֗T�H��)�Ȉ(N0u��7GQNy��>��y�/����pm���&��)����bw�$�$qȷ}�hֲ�x��js�����c�ݻ���4Mê�1m�ܜsO}�/?��|Z�H_;�{��EkW�9����u6ϥ>dg�7n|Н�`$l���T��1e���æ�rݤi��p��o4^�vUz�ex��B{L%D� �$q�f��H1B
� "�z��mq��6�G�ń��-D���AC�5*8k��c���<]|�����PT�._y���/����&��	o���<|EN]�И����*��d$֡ �B�����(��Ix0��z���Fk����2��`�(����VV�HӬSOJ�9],|�����є�ߴd֖�F0�.����f�u�>ȶI�-EE�s���R���˧�r=��tu���,��B��s8�R^��HJ���=PJSzYڨ���D�t$��l�1�,]�U�aU��Z�bzα<��=,
��p�J���$�2�@�8jP��؎"��I�9�Y&��2���P�7]&Ѫ���P���2M�\eQ���O�����    IDAT���Ԇ�BE�^�Q[��d�ݣ�h���!�-�s�����k���sOe�ɋ���Do>�˷�*y�u�����������]�IQ����E-�wz7�`]&�����~]V.�����KHIk8�M)!����	�]o=BJ��y���7���ܿ��/_�W^�ҕk�C�
�#�*��!!�Uak��d��考�Cd�:i=[ې�����8>>fuu��ܵ(�2b����Z����(X��I�0���9�Ej���H����[��j泄,��d_ꪤ2QST+�dY��/6~��T�Y��l<�hb�N�f�=�I����� �Y�G�*�:�?����tF�KA:<c����8PY��4Ր̽���3�_�-{�M��i�D�pT��NJk��u.\�ʅ�5�Iƃ�:�����fK�$Ǚ�f��g�%#"�2kA
A�
��閙���6#-���as(�&� X���K�q_�L��������\�P�����Wsw35�_��T�zEJ�k���8=;f<��i	;��%�=$&��F�L!���Llq�������e8��*\�K�
��z��(�uU�F�����Fߎh_��!MB3g��"c�R�&��_��s�h��$�H��_Wh��z9�i%ƾ� ��s�#��T��wl�*Ꝺ6�i|`��o8}���"6-o�M�GB�zs����(W�}���ZKD8x�o��ggԭ�e%#14Ik7J[����A����F4��$;^�������%��7�&R/J�+�TiL��{�0�r�F�F�	�˪�����j8xu����'��ƛ��h}��MRoÙ���b58������E��_����gj�k���sE���q�j��TDt8��CY�޽�_�1I�(�0 ��]���Ʉ"MS�J��Ņ�('g�{p�������aww��tJhjvv��7Xq�JY��'�X��O��h8::�6nݺ�b����:mF����6F��1}���Ί��<}�^��8ŤX��R���p���,+R�C]z�y���6k�5,b��?ˌMчˑR1���0����!�u]����x�99=b�\�\�h���^)kOU���h4aR�t�4��Q�'��WH�iGμ��6J\>Ƹ���>��Yk�rK�;��cLPW�D/��5!:GU��Fr���O�0*uS��y�&���ɹ���Ȓ²�9==��|I�-(AK�۩"dYF�4����K�}{�y6Zs���3X�D^"aP�Fw[qb#�"�C$��/�����|>���ʑ�%������R��鴏���$����1�k�HB���Ɛ���7�xc��Iz�I*� �@Q��k]�Ջ�U��a1G1��������O[����.i�����3�l�b��Nz�Q+����ELr�TB��E��X�{^�=�T�D�\�9˻�ڐ8B��>��!G�f +�x��o��?����ۿ�?���NE6u ���0���$����A�AU��9�I<��ݻ߾P��}-�LN��i�&�� 0b��(���0�M� mp�O�1��*:C����buI�n̼��X�sB�r)�wi0%�UD��-�FŚX.�X�	wr>������L&�f3��������H�h�4�r1g�8g�� ��Î�S���y�Z=ٻ�`�&��S���v1����]���C�`�4��q��}����/_����p��o��S�l������*�������w��DQ�u:�&b�a{{���{���?����px�"˱VX�k�Rb`�Z��Y�	��-f)u��Q�Ν�����VG�"�G5R�%*�&6�U�x:��+><���o0��&����������K��xL�˧}���N"��I�[5/�u�|4�mEȲ�,P9�3n��g~�Bb�Ν�L�...cs��f�Z`D��g���E���)�#vw����,��`�Y�
����`�� ks�/P��1_&�k-����] &�IOXH��*��ϵ�0s�>�<�=�z����8��2x!� ����E&[�lmj����`u���צ������z�]thX�}'ǚ���.=�>$bmR��\F/��ϡS万`��@�o"�vi��:��E3���];_v⾲y��V7u�s4u�K���S�����O�ۿɽ{��w�GY,E���9e]��#�|����;;ЄN^-I�9�R� e���pĨm�Vڬ�e���ֶ���_ݥ��I~j{�K�mmm1�88�K��0�Z-�:�A��՝|�Q�8�IفT�8	�ߔ��������m�?\��bϞ�5Fc��IPE��FU�����d}q��i��j��{?,T��cJO �����b�����|b�O��\-�,P]2���h\���2�,'�i�1�TAhj|]��e"X�����^F!E�5k��!fo���9��2�1|ݘ���y��H��6�(��qy��M�����> y��U���S>��C�5�Q�%��Q戡�)rG�Y|������c3�s9M8??������Z椴Ѡ--I�T'�:u�J�g	[�����1�0�&�'pn\akmH�s��6��1���S��Ӫi����݄�\�-�g��}dk���[��1r���w?z�Ç��u���� ��˳�^�&'��� ���򐲊�z�~rNc�����*ߪ��~�"��h����E���37�T=����>'��~��V����Sr�t�o3z9Z�QP]a�z���?���7�q�Ǿ����Z��^u�_�UU��kqy�G��>�{�d#v�n2۾�[o�`]��~��_qrz�[o����{+�R��I���J}�&����4Ep���R��)�g-�ṷ���2��s�dY����܄
�2�)�O���d��D6���,��C��*D�چ?�{��o_}�����}��Y��Aϐ���i"Ĩ���vn��:���U��u8�LY�E�J�YBS��K5m�.����^�ΰۊ5��MZ�t+-'�q�Ybh�c:�my�4z,I��� U"�敽�#��(�X!AlZ�s��鰜���fD�e�����ڶa3�U�b��5'ƥjHqX��E0Zy\"��N!rz��s���ɸH��1�!�����Ua<����$��hR��������YT�Ծ�	5j�@����l�ɇ�)�kmJ���{@c-�Cr؞ކ�޿���m�5���|�bQc�8�������F
5�"�$��S��)'G'���;����T�yn������	���&�-b��V+Bp6�(�LFc\fPm���Ū�,kn��:ǯ�����T8m�g�=JQ�֑e0�ʠ�;�*�r=m�^���������Ē��6�k���y�?�%�9���_e��ĸv´K�>����f��G�߯/-���I�Ŏ*�Q{1�/�s.�	-ԧ���tZP;y�""qMk4�VLg����������&U+��	�4MCY�}֤s�D��h�!/:�t�eh�����,F,��͕�o��:�ҝ��c�*���g-�Q��朝�%�WǛ�T�*A|1��h�yc�v9���GGx��}#�\�>1�bLH��h�4���u������������t��~�����j��N����z �1��)�D?�^h�bM��9�X��7�/���:�V�t�&�ۑ@;�в��g|F��q��k��"��k,�,�9����(OSG���]�G�<��6Q7t���Ʉ��m��xRP. ʍ�=�g��i|�3��nN��'�
ʺ��!�Fd�4�ȊU����prVS5���і3�f�,s��`]�E%�{n��i��^��N���t�~
-���g��^�|�^�=E�k�8g:�2�LZ'�����rNӔT�_'���l���=f�m���lIU՜��pq���R���D�!��4�r�����������X��Y�-��ç>z��iˡC��1v�i���4���9|O�0�����A�n�fi�2�}������`K�Mj������u��f�����Nx�i����K�/fݤ�j1�ĸ�uϲ�Xe�8$��$Bu����+.3�
��F�]�nȍ0�nq�`��I)z��ɰ�`�����6��7i;��Ј0�'};w�u�	x��|_�d	���9182;�����������{rxx���uT��i�U��\��D�ЪV�������1a_�wƞ��+K(\��[pѪS�(�����M���a<O��*:|"����%�*Gz��cl�N�`p�]H�U��~9�`�z]UM4�1U;~@Y�pN/��_�:g�q���'���w>��F��j@H���
�s�b��T>2��:�@Gm�e��J*.���`gk�ӣcV��q��֘���"����HSVI�c�3*�c�mHU��boo��(�ǣ��D9:>��	H����s����F�[�Qf[�:���u���dY{�����(�:�W���6a`��1W��l|�*���o���os��>��}��Pΰ�����;�ܿI����9��X��Y.眜�2�� ��l<b2as����a1_�������8:>e4�0�n���o�Z��֭���)׍��#�tU�=M�^��I�E�L���c#��'miQX/�X����:F��=à]_��+W�b6+�t��^/���c����\2B i|���`����j����A�n�~�����9��sv����C��n���K���9;;�В�'j�%�D���y��S���o3AI���x�����4M_`ש/ucbwm��L�˅�.���S���|ʃ���J�7����W�"j����y��7�J����1}"��N_�@�c�&��VET:2��e�(��һ�s��%�rլ�{��,6�;�iYόe8��n�?��4mg�!jr��t�i�:�����d��aV���_Ԇ�Ʈ��v�P.��e��y�q��E�����m+}2$"!�7��y�=�2�7�N4���<��s^y啄��}�|�5����8?9�p�î�|<��<�f�&����ck�1*�����4JR���l�b^��H&�c����2�Hd�loo3���&T�S̏s�z\g10m;��t?k�d� &�����c"pzzʧ�~ʍ�XqL�[��H��튐�U��PWy>�(<���V�"�!2�looc2a�UY�������>����nJ��bLh��q�i�ez#M�m3T,b��ω����˟�*R�FV�z��KP7h7һO�Fq��W����ٝWM�0x��� �@@/E��	������7M�#p��=�������������G4��r�r��^���s�>���N�_������HQ��������`B�������h����C��`��Y��������u����KwOuϠ�TU�0��+�DL�2޻q���%�M$��Tc�Ce$~*�֫�m_T�Jl*�,N_zG �[�jT-TԈؐ�k'�_�+һ_��=�#g"������Lb���iA������1��i���V�4����`Z�!��EZ�-�i$l+<����Cl;��s�i<�����0�ڞ�:Ƙc_Rvx]_�6a�ԆЦA5�DIn������GTָ�>�m�:ӟ�l6��A?�����W8#_R��0Z㌧Y�m����R�:��l�+�^��믃��?���^P�D�z|r�r���"��S�RMkgyb��s�a�x;��)n��9~�hf��ެ�E�,IJ'�iSD��'Y�UUE��d�`>_��_��������wf4��������8�Q�5�ɹ�w�����IJu`~v���G�D��Ŋ���G4��9��>�7�S:,T�Oc\b;��m`�b��^�]֞'�M��TXs�B?�4�}`�Tn�E����v�-o��"�_y�p��uI#>B�4�����e��@ދ�]�c�i����c.V+2W���~�F-gN�4�[5%#�|4�����ƍ�N[g�:N&#)-��#������>h"�6.��Y��ݏè�p��uR��Q��k){Ʋi��9F���};�Y�*ĸ2bVx]a`|�c
.^����;c�髍ё�ob�@FD4���}O���������s�����e[�aL�'��֮HumD�����������P�
=ۼD�>�m�vm��k��6gb/���0�������P�4���q�����4D|c͢�^�$ ��x��J&����{<M�e����9�W?�Ï>����������-vvvx���.W������!���Lfۨ"�\�|������Sמ��)}�^��1;�3�����6\RGY.�V���b���?�=.�$�!���u�,��t���	=�1����jU�8��jŗw��T%��2��5��[os���+|��(V�U?�؞mQd#&ň��4e���!�G'����Z��1�ęƦ�����W������v����Y�y�a���!�}��9{�J'":`���G5tYߒn��#�L�١|d�+�y�o�X�c>��'�(���N��F\{���ØV�CM��� &K�٘�2�/�X!�`4�����KCţ˰c>���.Ҽ.�3���1}�҆�	�����᲌�Y�Tvs����JU��>��\.�hGp�����39}۾�y�b�oauo��is��MY1N3�^�G2I��I�H�>���(O��^N�_��i�Ä́(�j��s@]=���YF>m��2�3���A�e��TU�)��G�Sƹ��(�\O�k"RU����]w�Wo�}��0v��h�����Rc���]�mM�*�q�MlFn�(7h\����qt�«#�r|P�
�qN�8����Ҁb��U���~�����U����|A�q�:6�9yh�����{_B11Gp�Lw���8qT͈�S��E�qc���?d<��ζ�|�޻���T��?���l���>O�ٚ�(k����(˒y]�}s�7f7���+|���|��g���<�����u������P�S�m�'_��ݏ���)u��{�����l�'���Ԉ����`" S�QĸD�'%�ɩM���9���޾�b^bl����P����)�{�67��g���/������?��r����9���|��f�n�����C&���~��� 	�b���Bye�&Lw0�Ġ��^��j�B�*�Dm5E�::������r{=-��I����Ϛ�j����^���a�4��t�|�
�[�/ɰhm��z����N� ������e7�=1�Ք8M�\r�6�Ԛ.sqUA1Q圭��O��l�E�N!\{���؀����Q��^i��
W�+B�&5��(+��?<Y�c���5�pb�pNaGԥ�.V�Te�J�d�f�pqv�a;֋Cʪ5�D�����m9�wo��G��[i���5�^����0�Ƭb�=Lt"��J`�R:�k8r �MD�W�� &�J'������*��)�#9E��m8| (HletB�rhq��I��E |�  ��vM8A��)nI�Gy֓z&,b@0D ��(1᪌ &i������t�0*����JN�>�ͷ朊}��w͆�䄏[߇]Z$qߥAŵ*[[[�����l6��4�����bӓ$�q��9�����e@r���{�������^����o����O(lRI0��j����N���M���/�h�hS|3��}?�N���_������6�޾�̓vv��~倽�'''|�ŗ	�8��n���::�)�^�L�4�#��B�A�}*ˈ`�
�v�=�ھ~�\�z9��}?|���~/;+�����q��5|i����-��>F%S�L�#b�)3�\,��ݴg'g�&�Q�h8#���D����3�` I��|҃+(H���Hh�Xc��Φ�G���9�˨����YKh&Wo�}v̀k�c�f��+�0��.5\.�]
$E�������FWfɚT�P�+�8�ڀq	�d�������,P��'N��4Q�t��N�a��x�R��� �Ι��ޣ��d�P�ȇ�����{�p��~+]癴�xu�`2\6�co͸u�^y�������{�����!�}�E��N
��d&�t��A�d�_�>:,n�/��۫R�y��4�b����=��o���%�A�    IDAT�G���p_WM>��3���|�rV�
I�Ay�X��Y҇c,J��'z��
^\��4MC�U����5a�|�_5x���=jCR���>+uyu����w�L������=iR2<����{�o�IOAT�(�QSˊ�k8�k�6�3;}���L'"���1���RŘˎP7x<�����FD#N��ƚ�K$4X�����W5�b���V5h��J���	K2_��^��^ds�VZ|��B�k��+�S�;B�QR䍎�?����l�����Z���@�^��f��"3�Pb�a�[vg�>��9��S�~�Ï_!�s'�A���I���X��>˲��t�R���;��w~����6�u�i�b�[Lc�m��@S�d�e������������*�5Tu�u��M��0}�M8�C�[z?�DIҜ�>6k-2��8�kO]�,�Kʲd:M����ϗw?㓏���Ç�:`M�1	C:_.����h4��H��D1��SʦS'H�^>j�V}t�9m��c�������t�ۢH��j�(��0E����U��{��l�yl����R�o8��!h1�%� ��K��|L���]�g����hM.Q� b�1�1��nVI¦ӇHO.��fEQ"F����$j�5cHd�⒟��ӈ�R���*�}�>� ݂t7_��&>f��!JΡ F����I_,�JJ��$�ISVT���D7@��`���|JrGѐecn����ɛo�f6��fNS��f�Gºk��~7��4�fg�~���rJ�k�,�h|�Ӕι6�k������.��$1��NP]y@�l����F#[d�A ��
[����N'hU�%�O�'F�?'���o��c$�L�d��9*�pZ$U�Z���>������!��Ox���s��O����9>�G�elMv��a$'�G,V�t����,<h��BL�Fg����X0$^�.�����3d��{�����[�Ӕ]�y��e{������w�.ߟ:p���w��o���Qc���(��]۟�=���C'Nѐa�c��D�-��qc�ߤ"O�{rz��qs�i��C�$��a4���
���k�T$K`n�o`�.W j���ҿ�H_��cΣ��7!`���S1��	m�"�fkUi��#bɊ��h��%,"4gyR/(Ya0�`3G�a���o��7�џ��;��Qk
g�)���y��6�B�v��"��6#˛i��:w���܍I������Z��f��k�1�N�Ӕ5>(��+O��XuT���sm1����6������՜�B�S�f������d�5��R��H�_�e����$|��]V����|���x��Œ�������������x�>xL���Y1����y���̗+���4��ڂ0�ku3�Dvxͧi�+qQ��k���cCxA��x�^^���Q���?��5���%e-�2�#}i���@B�^5�уj��\|u=ε���swf��(15��*�ڑ��Y���t�?顈��T��;ru4
�1�jػ�*?��@l��قH�1��󞾤�4��Z1<��?�B��.��jO�����)�ټd6�����t:m9���窍��F#f���,��w44�).7��#C>ʰy��##f�}�|L^�	V�
k���l+��%L�Ӷ���6ښuz�����ue���c %���)���0Ѧ<��x<5�!�f���c�������1Xê	��SV�4�4Բ��^{�O>���914D_�:6%��雉&��%ǯ�>�=��jQ�l��M$�����	��ǜ��p��=B�GI(�KV��*z���ǆ�ɩc��9�o��ݞ������֌����|yD�=�EL��Z'i:a�1M}KJ�?��H!׵}kl8����믻{��?d��i��{�/��C������F0֦j�����?�\�7i������5��	��Mcc���"y�H����PcA-!�{	�8�h�o�;;;�y�MN�/P2l>C�P�3�Ծ!4��b�`3�CV�)}d�'�4H��g�5�~i�1(���uZ�����>���7o�d2���j��0d�ш�(zps���(�F�J0IM!D�Q�씦ID�M�5���G��2�u�?�����-��:��o�=�I��K���ؤhQ��Ib��d�����K��%�u��Δ�*�Ϝ�]��#�9's��hރ8��
w���/>g>����a}|pz�G�9�[��B7�>���6i�fd�D�֭���K��9��6�"G5p��>����q1?f�8�i�w	P�b4X��Np��&x�:�Q��ط^g2������[�n����P-*�T�<K����a���tJ����k�k�6�k�ܣL�?Jm2|}Y��t���\��n���b���b�QT�d��z��������Y���{.�Ϙ�X��Q��s�w�i����T���*�4̐'���IڢVf��,�yU�3��u��9jr��r�����NL�80XG�ΐ��)RhI|^!HlSI!�F/��81}��;�.R8�MSr��^�Zˢ��b������7�`�X "�f��-��� �U���	wՈJ:m������A9�8g:��'��{����o~��X!�)��lE���z?���ͳt��H��g���MU'<��� �R�Mc�0M�}�6�Ir�:���rvv�x<f{k�FW��h+�8$��U��ǧ�/`<j鷼 �x��7h��DD�N�\�牠�T�Vz��*�:ùTT2������cDb�:���"����(eKW�qqq�h4b<��s��/EQ��̤ȹ�W4ՂW�~��C�����;�Ai��!���,F2��P��d9�h�+r����Oy�w����.�~��i�}��%3"��7��r� /2�s,�K��a2�є��o���8
/�P`���6�tL����<?/j/�\=�X�HUG����Yx�'�ߣJC�RH���M%Հ���!PU�шpnd.;5�90�F��;;�Z/.�*0~m��;��FM�S��1C���Q�*X�#M���d
��H(PM)L�9j"Zg�=֮1�A�s��Ⱦ;7UE}"��1@�$ǃ%D�
>�I�+O+ד�c ���4�Q�B�TƩj�e`2�$�SV&-Tc�em$%�������jj�1�&�z�'�|�/������є/;��4��}�l0}�u�M)6��o �������38=9O�![�rA"�jA^��.�����K���xe'��+�<�W����yxxLY�lo�r2��d��*l��A���/�ě�9S��bLd4cd>?#F�2��������4$gOk�@'�mLj��BĎ"�+AXGT%�@f�I�8=�9��t�<Z�8���ON��~��Dt��d��vm_�]�ܽ���ng���
���!�jko���bqq���HY���
92"��Ĉ+�;W~1s.o#Sk��r��}�D�w���b�QgBPT=���Gf���.� ��D�uf�1��)��TbhpbPIE ��!�>`2�8/��i�e��%��;�� �Tu@LҀ�@M�l�bO�>�+Fi�M�eY�R��c���8�O?������K/���8��g�/{��ED���{��#�n2�F����9��޽����z;�!yF5_B,g	U[l�f�����_����ې�T�"�	��TeHT%���t6�Xt����o*���y/׷=!�L���,K���HӔ�u�d��e���5����]mhؘ�����i�4��jA�@̦����]f-��kV��#՞�vm/�׷]U�1\�e�p;ϳ͞@�Y�X��1�A�TU}����ON��?{f�/�(6�m�bl#"�����L381D�k��✏>|���}k_.�W+��QbML��;�o�R�C̞�Da���e]�Tu/�m3�3��&���j��0T�Gu]3�����{���9���a��������g6���#b���]�}����\RUu]����O���S �˫�rw��� �qA�\�4�@�T,.��O�WDٮrD�d���>�z/�ʲl�w-���ޝq4>0�888�9��E*�0�~�~�!����[=�v}K��H����ΰZ����g���G��%w�~Ip��k��9::i��5M��*�
`�!�P.�|�f���<MN����d�x<���L�I]c��c$gwwc`U^�喦IrV1�)�l�Ř��X�\�ָ�F�awk�r� ����M���9a���).˒�bѷW792�	�k{{\�4�޽��⣿zO�>����yHS�g0VԊ1��)��{��w����z�c���=��W�FFmQ\�DH���N[�,I���L�,��pbhV�|�q���C>��"7�/K���'ڔ�M�����(�jY��S#X$Eq�U]᫚&�ӗK�UU���!�oW&�e�{��a4����*w��q�rY����o��EU���X$|�J�z��p���e�"�-ւ(�� !��^7�>ǫk�?�u�W�Ɠe������ۯR�%���#��Ƭ�ˏ��w�e~r��"bD��Lr�o�U��y�l��Eç��\R�O(�r~|ȯ�����X2�pn�b�"G��ܥs���4	g��"�o�m�c�t�у�Dk��L�,U]�\�S�Y�D�Xk�&G5j��E#B���qD�4U���A#�g��k)�N��f�v����k�8��ʲ�����qxm��U�c_�{gO�?o����~�b0F�5��&���n޼��ō�)ҟ�=��w�������)�-�<ʺl��1�5�%���5�bI��3?t<�x�o�ۭ"6��ǋG�9,��W���8ɋ�X��M]VU�Dz��\8�E�C�V+���\<M㙟�T��P55�npy�"�F�bZL`*� z�K��*��>Pi�f�RU�,�X��e�ȋ0��y,��Y�q)�g���dY�V�n��B�W�$����6�Ʉ���s��O9?����b�%��CįR��u�Z��zYQ5�De�8C%#����/>~���C��h��̦	b@µE-�l����}� ���Quiq�7�|�;�����cV�c���L��V%e�b<)���Q�d2�ڌ�+U��TR�dY�u�H$���
2��Z�=�1_��>p��.?��_��_������Š�9L�1�u�x5��ڮ�쉩�+
q������:&�K�cH�"W�5���S��oϞ�X��k��Z� �HTU���|�ѝL=b��G������:$3HV��Ħ�g0i��M�n��ih�y��o���%b��X���w sC���W`\DB�$s��ƈ� ���Ȃ4�4�@R�h5�h CTPb*&�*�T�8 �4uE��T�+`MFf�����p�����E#6kٸ��9HQ�<Ot:�ł�GGܿ���!�Zsc�(�E4]G�,����t9��H�o"M���fd.c����(9;:dw��l�x��t:�Ν׸��Ërp�6qB�b�6#����c���x�s�h�Ay��7�ۿ��|��'���s��U���kϲ\`,WgL�c�[3D�ղ�,=1���8'+F[$�-�Q^P�9���9��;����bvp��;�����Ǘ_|�~�#�#�f�Nߵ��ܷu�$L��w���'ڷ�1K�y#��c��2��o�[�N�ט�?{f��v�:�b���*�X��7:��|Sш¦�}І�dy�Ү��Z��XMU�Q#<j�t)�0Kǟe�d:����m��2w�0߾j[�+-�#�Z+�#��k��P<!`l�o�<y�J��u���I)
�!�DJ�V5�¤pX��@]�I�t�\���U�ˮ|�Ҹ]�9�}�z���)���dY���>�W4�N��P����9�t�Sa+w�Y>�19���h��d�l6�ƍ�e���)[�F������wU%�e����.Oc�Bh��=Ս1���͛7����;�&PW��Δ�����7g<.�
G��M)�-��	�%�fx��N��bB�;l+?hPʺag�s�/jƣ���h��rō��kQ�k�f쫜��c_Okݤ�Z����c�ƈ���Bhv�>���GnϮ��\�&�Fk��Թli�� ��4*D�Z��0��n
n�U��S 27�p��h9PhkNr�VI��AD%(fc�G{,�����X�i�@;�]a����nL��v��k�1�y5o�,����t��
:'�;��HL�A#�2�A".��?��Zub]�2�D��q3�����	�⮃��n;��x]{w�Q�z d�fL�H0�&V�|L'�r��9��.+�嗼�ڏ���f[�ᢺ��k�1�@�R��&E�@�b��''�l���MB��������bl8�4~������t:��{wy��O�h*��7�M�Z�@�'9����>� d�\��_-ɳ1�2�8�|�v~l��y�f#���!8�h*"ڻ���N"���=`���c2��뺯�"�7����2��Z|��0����ވ�Ez��L�#���YY�U8kɍ�=���>��|�/��ⵢ��:,[z�W��1�JQ3������ʠ�x4cȓhyb.,�^�~{�=ɋn�	��(O�����/ُ# �t����ߴO�� R�} 3Bp���E`���Q��&XS�e��UxW����?�y�{��5��OĞ���{S䙫�1*>Zc��[b#q-���UX�a�eh�^v������.��[*i�H���ገQ0���V�&��ld�1;Ƣ^9�H��!�n;,���E����988`6�Q�k��,���L��~�mn޼�;�ï�ׯ���ҴE�`ggg�6�,�ma�e4�A"�/IIB1��\I<b4U���k�:M�}�1B�5>4L�#|�F��������`2���$��U��Q�o,1
D�c�T�h�(��`\�ƫFa2%�ؤIAfZ̆���hDY�,�ˁ��z���i��4Mr>��#�Yv������o2��uXG9�e9�*B����},Յp���gv��E���K2.�2hC ?j	��ݴaz���u��/�Jr��].�����I�52t\$����!JE�%�����?g�H���h���Ísꎣi�6ř����-N�N��S7%M�B`kkь�?��w�}����_n�\��'PV�1�,3��cb�+���Bւ���K��ڳ�͋("�!�,��|�޻�f3�g�̶o0��߿��=��%U��E�t��6�x����o/��yJKR뀸Q�~z��,k�j���Q�1��.)˚����_��8=;&9Ǯ'��a���x��]!O*���Zi���x�i �<C�Xk]�qbȂr�!F~�_�������OĞ��3��7�I"�1���E�T��=�${����m�B�N�l�L�pi/n���f}�YqI���rT"Q"Q�zNY/�}�ƒ��SV��ƹ���h��|� �EU�V�jA�G�N�Y.�NJ�+֦������"b�1pcg�<��f�X���i<(�3v�ʀ�a4v���INP�K|(���
Vobrh�}/��M���O@TT�s_���rt|�'}���vw�x��g��z$ɲ;��9�^[|��-2kk6YlvOw�C�%B"��a ��[�#�A����y P�<$j��iABJ�fi�Iq��j��fuwUu-��ofv�=Gf����UDdFd�/��%=�����=�,���ob����loo��u��޽��l����x�Z�qU�ށ\��h�����֢1fޖ��*E�r���>{��t�<O��!�������-�d]:��xɕ�=ǵN"�u�:bb��u<�����t��2�܎Sd��I �@4��j�U=��dǵg�*��tQ�Fg��f�?�"@Ϟ=�t6�phaB>L�� ���SXAVa���H]U� �AQL��_$�'*��s1���Q�ʢ�?Z� I-zY��J�O�0@N�1B�D�"v�	���w�q����CiP-k� h�	�z�]0��5��@9�FS(����� "`w�)>��
U��ܹ���h4�[�-�R�4�p8��=�y���~}~��ԲIm;�v��j���i�����柟eOD�    IDATB���rV���^
k�n����BT�bTUk�s�5�P
���lx��A���Y������ z  2��Pa,�)�O��	x$����&��d콟W#��*w�2����X�9P�
Fl��	9!����e	@��C�Z�n�����F;�L�_�V����PI��=,�1�e)����
�H8���3T3f��k*(��H���D���~��;����7�	�����!�=|���;��U�髯��誥����4 M�
�bŬB�B1��5��0������a�;��$�F�3uol� !�ab	A�6�k�I�=��pi��u��Z�� e$V�������1�.��s�6��x��9��)� ��|�s���e�䝄��'Q
@��a��"�"�,S��͛W��v���W�z/!8%�* D���(����m��������
ۖ�*�8Lq��w���һqR#Ԇ>�b�<ϑe(|T�߸��~�����;��t4; ��\=<�H���$I��iӓ�����|.�=�L��o�7n��H����^�\�=�=���;�ֻ����|@ݲ�52$��X�D�u�PS�x�������b�B|�?�s����B����y�$"F�H���3(	�� �`!^�� �����E�S���ܓjc��U����	Q��!��7� �Z���Q�T�^�7n��t:�{�F��"��hpG�kD+aԎqQ���2�<��n���d���~`�k�錾�z�*U��V�B�D�(s��{�XΫ[�������úz��W�p+颵D��AF��`r�JE�;�o�w����.b9Äj#�(j� I�y�d�=vvv�OZ��s�!�j	�,���E== �L&��X[[C�� �3��>���.{I�!1)����d
�dpFPU� ��B����AljA�3���*�:��	����g���� ��>G����p�]�k�
H��
��U���A~��c ���4��i{~�6��Dh�Pfn:�� � iB���I[lT5������1F|��g��f�y�fc����u��\�H�q�ڕ�"9Q�(��T�bϕ�1��_��\9���'�1�5�� �����g�U�HI�`�=�u�I3�:|���"�<:�+�$I%Yr���4�줉ʫ
-΃�>ŋ��X��D �ß�uv�"���XW�Ɗp�7���W��7�o�c�����7Z�+�v���4=�Z��m�/�~��q�1l�s�w}�[JD��p�U�M���d2�͛�P`2.����|���
����A�A]#r�Ź�q���n��|���`!�����)�ky�Eч6�#Me1ڟtt!w� � �}����X��펡	o��%�(s�&4���RK�4�i�@u��$I���������N��أy��a���뻼�Yu}~.ڨ���q��w�ߟ5�q�y��H<��,?�X�Ԍ��M V�9��9�z=$���g���!�4�T�4}eP\]���������������w��>@������.�{�ۿO��v��kU���p,�u$t]����q��[���)qD����S3�xv0b�x|S��vt�\�
!>/.�-b��x���,��v�B��ԤU�DX��a�����h�V���b|_Ǹ����o��Eh`�~�Wu��A��w�Qp�kG,���i,����݊Dn������PE28*A����=�TM;2s���|Z�r�Q����K
��*n�婳[e4.m�1�)���&|׺H�̊[[�uo��s,���풂��L���cgf�S��f�Zs���O?@٦��n�´��@���wtA�3?����i0�3�f1��)�L����N�
��x.61�� �C��$�a�۽`�K�Y!����D�Y��8�p�Ԫ�@�>t��Պ4��Zԅ��5�.Q�������;�����q�V⊄��ەK��g�R�4��o~� mf�ciߗ�3��`8�������sW����g�$�~y.$�Dishq#�ڻZz�P6����?��iM^'��>U�)�������VK�>����Ͼs�G銼�d�+y���n|J�k���|<fn% �"������ ��
�K|���WB�q(����"Y��e-�hM��Sm5w��@1w�&���%�>�q(N�_,�ڗs���^m�_�1d��F�Y� hjd̞E6F�����E�<�K���R�İT����eK?�t�*�r���)��w�X�m�&B�d�5#2}����ü/�m�ZZ)�>���35�_�֮�9����Oj�2'K�Y1	ͨ���Y����c����u����U۽�jl��܁��|'\C�UDJ���DpD(b�/���[�����q ~�HJ�_�I�6H&jjf�p�dBI-S�q��*�l�H8�����ڍL��H#p���o�OX^M�x��4V4�_'*tvWI�"�Y-hXT��"���?�&�]w�ͿMb���չ�+�C� � ���۝&�m62Q��wd|g�����Z�jL��͛�$�q���J9�eV�����d��{*a�bЁ�O�e����l�2{�bu��2�P;�z�݌a����ݿ���q�m�SH��� �n�C[���f�F�Jg���h4���*�𱱣�Ш�H��	��U�;A�0�c��W�B�������MqX�մ��!���D?*m�0�`�`YMa$E��g=� ���9:���W-�%��%�����1����6�+��L�W�%jf/Vu�0�u���s*��
��
�w5�F���v�e=����{Y�수��,�5*a_�j����*�j*lU[��P+,س鴪�9��y�?^��p�Z��>f �E\�r�"��Xq(�Z�k��}e>��Bɮ�V:�k���T�"E���8M%�M:E�i�􅲯B�ǰ�*=�Z��O���Hl8"��� \V��:%.y�����t�Z��_�g���V>/��W'��9�C�����Sc:�.��O�_��������ާ�9�ִO�_ZiѸ�	!ı�h��_��\�?���Y��I��W��G��}�e�h���[�������b�lQ��o����R&���E���Y��u��;�#/F4O&�7J|LݽD�:��\U3*]f����0�*�W���P��*���}��{ c�X%|��P n��1T�W����k{��֓��|�?*�{�Z[lO��k{�׿1�g�%��
�+Z�_,�Ԥ�Z� ���^I)k��g��(y:kƭ�N�ؠ�O]�j��j��HK�GөzGǗ�������B�X90����܁w���`{i&a,+;f>j�h����d'��%W�Qk��9�L�W�' Ai�gq�F� ͧ%�����f�u�o9.��)A�ny�_��<l��w(Y��4}A�^���h��ύ�6�"��`.��~یl�Kk�D:ퟤ���5q��l�e�:pF�� i;.�A��/�3�SEu�*5�^���5cC��~dO�^��S��#����֒$"�*�qP�7�o������yW���WM?��o�rMcu>�tJ��.-����x>dp��|���?�Ό�z�fَ��9p�+�̓��DPή=mO�����\�7	�FF��M�Ց�Tf{��RKE��:Z����<{k�����o�{{�B{.���vߞqU	�in�P190!΢miL-�O9j�a7h����1�}��z&L1�IF�)V�#�)����!��4v�Y�Wn�P#��P���%���.(���VCϕ�J6�=�T�%d�*�+�f����e�=k��Kj��צ.�92�6����
���a9�d����Cz2.�@^�QoP����)P�<+'��xE�'��=Md�;.K�E���x���l�HEt��p�!��O34"�:΀7M�sqlD������y���d�XN+�I��%�u�<�qve$q�RRi�/��4�ģ�o��XkF	�E56R`Vh�+d�K�-�t�s�S�6���mK������jE<r˳���C�,���\��P�Ilf�;�. ��g�zo,�eTE3"7��Q�Zьm��n�����P!P���a׶��G��3�B&��rK\������}�������GF#�����{\��V�D�Zp�/+m_E�[X���Xִd>��,��8呹	��l�K95�~���ңV��sqC-�H��fh�~����C��r-�����̕H.js6��S>[;��"�(hmB��%<�M��u���+D>����
�=�Ѐ�˱���,�����0� �o��D�	X���}+�$IIIk8�SW>0{X�%����_���˷M[ �}��S9�&S�I�������9�����sN���|��*!�4b�a���L=_9^��$��ys��q��b/( ^�և�>��d;�����d�E�T{V��Q=�r:��l"�Ft[Ă������9��Tg��/�����'����!�Yt����!�YMG2����p�´[���QDJ�AM|J^�1o�}�ƃ| 1'�!�7��G�7|/�X�C$L/��j?F~��ώ�'�IY�gã�R�"�d�d�ꆠ�:Z�ĝL��?�}zS�ëq� X���λ�VZ>-�g��Op}�S<��	Ƚ��611�LB-�K��v7}��탿��1�qq#�۝��]��*y�rF1Dg̽%�ʲ|�Tj�@����z�\
�~z��66$@Ʊ�DՒG�_(SB�d\�`2c�.0�=|f߳����W�^�j��[L��#g�"���t+�X0���˚� A��3u��L���|�j����C!�&�t�D>,�Z�t�������)��I=��C@��ǥ;��5�}:�}�[�h��B�.2�.�AR�y�!n�.��.\�X!=g2�8+�ThO�Rj�:�¢1k(0<���B���E�H��2�!-%BχŀZ�S�h�W�>�Y9��_���$�i��o,�=L�y�Il� m��8d=F@'�|HR�`	9��P��{��8�srѥd��t���\�ċ�� ~X��ݝ�3˔0�-�͘/�J��O����x��ƴ]��[_��G���v�t!lUP�I�2�u�/D Ք���L��(E�LG�7����bZ�\���ȴW5�,�\[pر����qد.���y��O���f?l�o=�~E���}�F�����>)�uS�e�>�����sڨ:TH�_��m����E�$:i�]~Ft�zҸ��p6a�I���Z���:u_��,����h	�A~sbR�U���~9o��E�uN�g�������&��d$R�4E+�9R���Xȇ$�/��W[�^wMY ���DY��aG�}~�����}̓�>Қ��o�tn��'6�.��`q@��4�@t����<��J�f�rMو�����1 e����Y|���z��{7�옾�Z�o�����:G~jK�6����TM���f������f�LF@�D&lX�j�1�3��Q��NJc��+1
�EL(�Xj�4���_l��C2H�-v.�������x(6���N� CJ� �\0�Y~j*����v��`�n�����3NRlWR-����������T������Ժ���WeP�DH����$۵��K7]�h���9�5۠�܊�����i��[/��.?�S�0���j�~a�FY�	<�Y�kGƠ�?��+5��@|��`�ge��`,VN9�3���$O����_�����q�Q��0I��Y�_&R'��K�>zF�
Y�T��i`G=�ĥ\�`����~�x�Yd��i]e��� vB*5�$;ﻩ����\��$\a\�� ��4g�Rj�V��\#�%%�@��|�P#)��q������8�W-����q�p$,�"����%�$�/�#w�Q�!���>���G���ĕ�C�~��'� ��޴#�&p� �zg���S#\e���!
��s:۱Hi���DT2R�������0��1���0d���ԋ5|e�2tvn����������������d����L��Z��2��1nf��CK�hp�f	;$�K��^�W�9VQ�1��r�u3�u�;��S��(&��	je��A��/_��Ӗ�Ц;�eP��U�[��b�A�d���1�����5	<��g-ԕ ����_�x�&���&hu�чe��]Ģ�?즽w��:�����]!� ��7�֎g��wGPe�M�����8��׬>��f�P��G��(����Z��k0�_��Lw�����'��w������ܸ
�gh��sUceLM�f�M�5G�g��ݙ3=�!���Rm��v�K�׿V���%~0�VPQ������P1��f^�,��� $hf����,{MkۂA�?B�y�X5�9׆�T^��}���SAy!c��Ie�������,��K'�6LY��2�z�+��Eمϟ��Ѿ��<	Q�����A8�1'�+��j{h������2��K���C_�(:o����������=,~���X�o�/i��~��ۧ��sW�a�`�@��M�qF�u'+)郎J��	��n�;l�Q������7��P{�:�H�-�Le�]���?����zo���@#����x����X���GM�4+����99��PX3O]���P|�Z
V&�n�e��Hӵ������.�ҡ�`E0+�i��0�}hq�.�
������0�L���n���/󾦫Kv��]��;���c���ZON����ޘ�������)�Sa�S������O��8s����_��/��������D&��v�[��v��{���|e!HN�vWx��3�P�lwq}�v5��V�N���-�T1����7�w���SߚF��{[%�̰x'B,^�G���N��UZ �����A��q���^��
�)�Y�6���Ͻ� [�������zݰ��	t0�QP$�W�l�lu�W������f(�)�Oo,>E�!I�����!��g�bH=2+ǚ׳�Jg���sC�e��0�)G��2����� ��6K�ڭ�P��;���@�2��%���p���~9��?tn7�Z����m4q��ˇi�\F���PzׯT|�\�J����K ���p^�H��͕����t��Yā>�qk��d�K��&SX���Я5����
��x>ێN���3�!
�Iy��oA�M>A!���:_L�w��}��8���H'�
r��=T��U��B9#)o���:��'>�;�)������z��Ҥ��!ɆA;K�WT~V� �VӀ��u奔T�[PwY\���ڏ73���A8,������i�!>?��r����n��g��̼Y�� ���qbuZ%���4�){�?T�@gQ�4|¿ո��`���c[V��4���i�s�������o��/�,�WN3��C���F8#(�l)�*��U��_u�5nZ��o�c�Du�&�[�z��O�/���}ă�ݏ�}y�>�?����u.ՕR,�1���N��Mν� .n�SqG���d�(�M�$����#^���<<A���͇��n��M������$�����x),����"L$�V�g���&�Uj�؋@N�U����������܌H�s�/����\�E�����moΞ�˓��:xm�WG�83���Y|�H����;M�:JU��r3Ҙ&�@$��Ÿ�y�a����2�:�4����%Ȓ-� ����tb�00��
�+��!�ib@���{i����ܬ�,H͇�j;XM���I5�?����@�tq0�U��Nx��i䕿g;'f������;�&/�֫Yx��DG5�t�I�p�;������e��"l�}�]�b|[O*|2��&׬Xo�"d�H-�����o[\YBv�|�o�7,�(�sh#2�T~�ڎ���3Ko��,�IH	cr�C=\n̩h4����Dگ�x�����-�'�"���k_�ٽ���"S�k�zW�6��ab۵����fK.�I-o���X7�)ŷ����U�-��Z>�v�|M7Fh(�U��tj\ﳒA!be�APt{�/~x��Av���=�^�X���XL,DG�'���G6�8q-�̧����@�m�0y�^K��������EG�uM�~����w�3a%�������ƛ������LO�g��n���n@*'�Sv�V�I8�]���.&NǞ���ã"��/��ؐQ$$k��s���c/���(x��J�յ�Ⱋz3l�G�RO�j�Wb�(�#��X���%A����o�&��s�b�>Z/�.�h�_��W�g�Gy哒!a0�R����7�g ���� �0�@�,�n�"tg���������)�+��5r<T#��ߔXɵ)0?Bo�F^�-�`0<�@�a1b���ƣ���i�D�#>g�1-�膷��j���.$�-4�����}�Á��{��Y��N���[kC9�퓓�	gj��FZztZ쌼���2����G��̗���\l_ϣ�߷��'d���Dh��m��0M��T}�5�#J*i�J�w��Yp�%����k�5��9^\�O��U�rt����rKK޹�Pm���&<�(v��+t�2<cJ�Oƴ}���9fg������4��j���ʚu$nG�
��џ�O���u�aJ��
��v+�O�GQ�����TVU-H��)d��֤��*�n���̳k�*�T�Z���.�5�x#E�4�c���L���I�|�*�/[H���C��G���^�*H�'ͻ���U�)LC��iz�q1C��o=�e�o�}2y|�3=�M��U�QT�����ݲ�L7��\M=�zmXw�c�I;Vj�P^4��e�3�S��/�Ic��`:���_���h�~sq������u�ϲ3/����v�<�?�NED�+?Zߌ�s �N+D�I��(�wPD��-+�$|	Y�g�$6+��.?�Z����t�3`��<h�Fru�E�K�qÚK{w鞭v��
xF�v	���"���P�D��pJ�Е鉜i�r��g��&��Ʌ������pe����'�w1�A�X�JAV8 ��4̬�����O5��_�89�?P���w�c(��f*�3��^I^���L�{M���
ΜO����n��oϪ�c��^��Om�?[we�v�6�������3r�w�\���l�}F����z��׿��_6,�����oq��-N�O��	���&j�S�\�Q��N[��X�j�xवc�<|���UИg���]=Y�s��`Bx�56���l;n��κ\�9��d}�/�'8 z��MNO����k���$B��u�qiC@��%����1)�F�~M���A�����@�����`z_Cn;]�wI·��?I�`\7�������E����d��gK�����1;TnG��r<���J���H��Ժ���y׽��j{�H��(Cfd���o�K���;^��9M�@�CS�����>�~n�q�����S蔒2&V���1���^�e�H׍rĵ`^����M��1�������z��E@Δ�-/0c��d�P�7EM�����w\\�h���&�����g�@{�ȧ�5�}����:��4��Sf����f�.�+�(�X~�/	��_�Ǆ��lJ'Q�4��18±<��+�_���	��<H���qo#����?MŃ۟!��7G�ɟn����ݽu��	"��m�cO���[�!/|�����6�;�
������y-��T�v���z7�ĳ�;��G��CPx(`�*!��yY~e>B��	��l�����{�H�@Ҽm���r�'n>�;nő����0"�F,��@��򗑨�Xh����Q�T�kZ�f�Q�Ol�����I@ȃھ���$�{� Ʒb�n�M;;��@���xOk�3����z ��o:��u�a�O��1��d�1gk��v�J���|���2�  hen��86�sJ}"\[.�+sL���}]�T���$J�+�3\:S����{�*�	z"�8�|fA�2K��.��긶����ո�3�M��5�e�x�|OƝ$K9Q���.J���F�6��6®0�>�
�؏ �{Q����q�oh���!M��2�'y��t ��V���Zy������򢍛����Vv��L�� �{.�3�7��� g�1y|��|g+W
7��	���xh*�s��0���T�w}� (rm��ӏ�b��")��k����JT��p	�H�����8 S�9Z'��B� �j>�DCN��J�#Lp�HlS�$*�D�'i�� ���#q	�$��W��G�ogfE��w�t=���yI���dbb�DS�c��9g�˰��n9޷c%����fb�(�w��\9����n؛��s��zF(LV�.}r���^��^�n{��vݴTX��jB��P�gee�e�@My�m;�ω���)��xy %�������)}�JO��?e�`ᡰz�,�D�VZU���o�Nd~e7��F�V��	�./j��ܲw�W�դ�����񅄈k|�*bb�+\T?�˟@E)�\y��h1�EB��'ؾ|Y{ۓ A���Ɠ���wϽ2�F{����aƶ��iɘtm�E���s_�&�_�A5/[������o�h��hp��ϹJ\S���7�";���ʡ�ӝL����ʙT�����L6R�I��r���l�?bA[̘gY�
Y�7@=s�P��Dl��ׇZ��W���K��!�=2�&1��G��6����h(�?��\�c+��R*9��)#�H YU��y���>��E_;���  ��f�j�e���Yョ�ޡt�x�_=|�r�b�
�7���T|'����G�
8�E�,^-��\����
.n�ӷ�5�A���z_!zSO�宩�f�I'":��������H*S� 0E���?�}��E��_?�U���7�W/�Vqf,b��L�4є`	M"�/,|n��	�/**��f�ṷ}w=��,�+fS����ᗛ���K1��"B	�ݎ��5Yw0��L'����:���k���`ᯮ6�4�W�s��X^��Nط�ѥ�^T��vPSp�<� ��iU%�����g�MFu��4��]cg�-���iZ`�K�B8h��`�����u�&CJ��a�q���x���b�q�$�F��]QE���F�A��T�́��2��F��F{��i��l���/}�H�&x�@+0i���s5(�us2?3r��@F�B(G�o�=Ώ��E*��'���Q��SǷ	�����Z(�X#�"6����y����S�IE~J*ݤk�O�t&0w.��O���(ͱ��0��6W.�A>�����J&��lM�6[v\\_{up��F&�A��@��ꭞ�,#�M�� �W���e������c���Ǥ���3�H��j��Bz���NҬ��v߾g?�:�N�l�W�U.���jp�59���
QMѶ��*�%��x�cn�u���"j�<L���гhtY�w*��$*�B�Ԑ�RiԬ�(x���hh(���vu��͏���rۀ�|��_���%�<V�JI�L��7_|O6s����mЗ��;1L���������㿖�{t�>�,5��?D	�{��Y�E����RM��� 5 ��܍�E&��M���UC�!j���d_z�_����ƣ��`d/�\ݭ�_7�v�q*���Yt��C=ӌ~w<Ɵa٣5��5!3�Dj�A�J⧃͢�5��8ס���yՓ�X�$$Tl��#"��r
�?v��5=�c��0� 0��!�"�ՖI���í��)FS�&#��CC���YR�r��-������H�\!�r�9�+|W;���h�2�j�^���ү�̨55S3��x2!�y>f�B�~�@�A2�,���0"�h��	�����IB��@Q�v]�rGH5��eZ٤�5�����\�����E[���2�j�|�A�k�R˰k��0u�3�A*�r��}����+�߁���3m�-���_�OW6t�����7lR\6�gw
b�q2�tJn�]*�X�G��;��=<R��~:;s��q��D@�8h_��10��1��y�Vl��.Q^ۖ/���uo��s��מ��T	��xV53c��)x�e�W�V��A�� �j;�[�h�7�(xo����5LEVk;��u�}�����<���HI�
�Ї�^�@xq�C��d��8/K��*q��=L�pkqk��g��g�Bo�C�k�B���Y���G�����/3D�\��v��}�cTs�"�my52�M�@�T����Ǽ�܁-�ʋdݐ����=2��v	?x��g%�ӯ�_�\�5��#��gU�j)�ȋA(�yS�g�l* !_�]H� �i��S�qs�,��Od������e-�;cFY����'�2�j�޾w�x���7��\騿��ԁ���V?�.n\�s�Z	MJ������5�I����>8��B���w����7��IOg�O�pG+���A��J�U�I����`*!��'�G��Y�p�0[�[G�*˅�}������4���1���N{����
_�Q�q�`�V����"U`*��g���wm�����o<�nٱ/in�&{���_P���&�Ʈ��P"��bg��(xڔ�B\FU�s�m~�����n���I�'��n��|��#U�<�>��T�-K�3��Д������SB
��<����2-����Z.���0cY�hZ��7�m[���X�K����͐�iu��铍$~Ԥ�Q���衆�M�S	(Dܾ^޶6�0U�^%�����'���n�=�0=N�l��T��\L���$l�����bM^<��ʥ_�#@!��&�(���8[�ވ;��PV:�1}�Ye"��K.�Sx�8=��
�<��tC���4��İ�j�$�B�|��	}u,A�����O��mc�B�T]��;s��$8(e��Z��j?d�q��6ӌp�#��\1?`l�^#��yÅd��Q�ح��Q��R)�g<M�@�ϵ(y�����s7�N&�q-jY�~e*�,@!
�*"$�I!�/�z5D9���f�ņ�l�Ww���68jڝ��0�K����*�Y5�O㨕*{�� -<�&��dX�^fs�:�Q�����_��&Fe�fğ�J��ۺ�I+�rp�^�܉�s=e;G�����`.�
w����J��q͵:t,l�P9�>-ڄ��	����7y�o"L�j[:���ow�s�\������HR����K�#&�K`N![^�C��LȘ��,؀v�%2$7>U5�������d��gP����Uu�6aF��J^� u18�����^�uTDxX�b�/�U}y(� ��uh�.��if��J��1P�T	��CG�ۤ�����*���M�%�Df10��E�����l��d#���5�������
c{�<5zW	����Z۝�iB�#�X�H���	--���|�����a���0o{�$SYm�kk��Jo�%�����
��Ad1�d'�{ƿ��g�L�����}�@���	 ����P\��pȎ�k�Nmuz�|��N���wnd�l�5��-���D0�%�L �T$�J
1F�%�����&���mGx �ƚ�հ*TJ��a��%?��SW	��檜�Y���3�!=�^�_����9�Ʀ�R/ɊO�vU�v��Y���K�߰Ʊ����E?iW����֠�%S�%P��Qa2����#a���#��uA����_���[�{{�Y���I�Gc�0p��۵�KX�嘼1�j����M�n��rYrl�����C�� iZ�*�o"��s3Ɯ����C]�������Y.�����=~��������h��h}���P���r���&>B���D�A�?ov=� &r
�o�!=(s|�g���,���ɀ)��A�jր���xr�Kޗr�!����~�u2�-˘�����y��g��66S�>jq���SaIY� (��:%m۪ʔJR�G9�X$b�ԩ~�K�Z`���[*<���W�D�-j
���^vĆ�!��>o�Jph�Ḛ`@��,H}��@�?��9E@'����g�+���HMU�.�)�5c����hC�<:ں�b߽i"��q��3\�h�����{��Ǖ���#�� \�~ؐ��U���zv�V��~�A�{�_w��NrM��&C~gn�C+Q���b�)[1�HD�G�G�΂���0���c{[ۢ��m�X��Ȏ҅��bP �Hi�Sy
�;9��"�W~�	S�
���m������A+j����sL��}\��D������{k5 yxx�&�?��o0���ݧsl�X��
���&Ao� �Y����7���:���,��M:*���פ�Gs��GA~f�Fm�1^'�42��yq����d��Θ k����5������[��,資�&FfZ[�=]Y�X�*�=#�r]�5pM����-�y�嘟�������w[���ލ?Å�I�>��(�hJi���3�+EjU�ɨ���'J��%uѦ��Z空�����n���eu/-{�դ#�5q���7��w�/,.fD3�`P(E@�����ݽ���3��_מ��k?;1���VW�2�ĕI~�p�2EAO�~2	od�?���'��N�+��܆r2�48 �~� A�%H��1��1�L��T�֗a4q��~�r�v|�o��4!T�tU��GP˛1_�؞ߞ�w3U���ԣ穀<Ec�"��/	���P���al�T4E�����ݴ���ܘ�5�1Y��+!z�:���ɋ&:/42)�����V��3�t�Tj�*.O�F�\M��À��*���L��K�*�w&�	�[l��H�����7���W(�B��?ц����X�w+�y��#�)O���GQ�>MSCq|��GI����M���뭨;)Щc�E�	��j��[7�Vo����	��ʯ�{w���b�C,�l��E�����@�3��j�-X�~��_����!��r���3Wq:�wI��7���Ns�|I��^�}�dO����$8�r��v�̊�H���p�c��7��O�+,��Z�;����y�7LN$�K*��IHF5��|�@<?�O@�8��o�g��z f�6
�����'.���/S�Ô�l����<���;ã2����,£Eb1f�V`��T����7�)�7�2vL���+��ŏ �������xu��@���w.�`F��<�$�#�h�:U�&����M O��T�Ğ=#�̫H�LE1SI�k_���}>���H���=�g݇�u:�ɔ�
���}���,���w����B�ϻP�I�*d�y�\qX�^���to�q3�a��`{�%���z}���sWmt C4T�OT50=LR��-�\Ǐ����ͩG�?�#�J�ɦZ5A0�t��F������y4)`p��*Ԅ��{?]Yˬ���W���ge�T{�uv��g����t9����˄�5:�A�^�=�(t��beK�4�l����u�6�j�ءL@������eU*S���vX����d����OjS�S3�L�0�:O��"��=w/9���~6�CJ˭�Ic��o�`z��{ϡ�M���g�vE9���wX�1�M�!̮Pm^ٞ����L&��"c�"�t]B�j%{h�����Y"qlG�@"���o���e�Q�b%!!!FM��D/�)�9���(=�/p���+ ���ږX 4`�?�����e�g�\�i��+S�k�u����;�`�.��Awl�D�`|L�Щ5�
طBƙ;G�׾g��G�c
x7?@.�Ն�~���h:����KjKYI�/	ɠ�H��H��S�҉��d��Mj��9��
��v�Cw�JQj��w-?�ne�=U�3T��nF�	>	���@q�M�b�*�_��<GlO��>����R��iQ�6���?�N�|_����9��顦 ����R�*(�f@���Qڿ��6�έpc��D�:L|�o�P�6�|�{-�y#;��Mi�3Noyx������k�8���$��ּꜯ�w���k���B	1�#Bm	��qp�t`�e�P1d��v�P��5��	�٧z��Y�)X*��bD�|5�����3��gS����j�Xb�z29���Z����"A�����7^!��M-J���1u���4q7����&&vo��W���~,&1߇ q�u�l���ۗ'-�]_�RF���Y����H������{	��3���]�yp��lk��g�3��$�[O���OJ�w���k��x&3��q�H�,At �`�a!Fb�[J���z��ũ	|:@4G��9�OR��0΀��Ҥe,&�8s��C��^��;��@ׇ�,���D��I��@=�Yo�q�۽��ΐ��`(�sG�{��նVϗhv#u��6�.�S����sU��^��X�}�!�I�O�Ԕb$� e��YKz?�̭E�c��?妥�E"6�� @��s��%=
����#p.�� �X��ئ��\P�aE �!����]���;�i5�m�e*�������Hi�P����b�3؟iV#�ts'��7�UظѮB6��lK�����y�M҉��j�Po�������������g�r:��f��8H�H�C)5]�����z\Cߦ��*/TvD�H�V	� ���&o�������?�Q$n�5�Q0��땢�
W�o�99�[7&��`������M_�
wy]#i��}2����v��PZ�b/^�ݙt�����yt�`$��*sS8���z|��I1Q2Z��Z�VG �y����vX,#R���fX �B�ŤX�X�?�	���x�:���N������p㕈HA	��iw�d��t�
���u����_�\4�������^�	?�
�M�e�~�₎�a�ο�	��r#���?��x���x{{k%����:WDi�\����_E���5S�U�YI���/��7�L?F�8x�7t��id�Kf��]X�{�W�|#�w��Տ���B�աINT��ֳ�}�22!�Lma���~x��7�]>O|.�S�`��7_�?�?�5�z523���7VG���]dޅg����$��c���5��p�Q� ����C�a��~�i%h"���u՘�-f�z}���i� �����N�;�z�r�Է�pD� t<�8���XI��:��)��P'�	
#��F��J.�<n�FO�LN��bݢL��A�̿ ����G�Z�,U�����	�G�w��$�"�EO�C7��{3@�ۄ=%y��&��lۗ*����؎�%��]S��+c`�N�hy/�Q�?���mCٗ�)�C�&q_{�����[l��з���J)�H�d�ym�ˊ�(�
��\�&����N�)p��z_��V��~r��	�}���b4x����'J��I)�)���O#��$�\��=�m�����������m޶2I|��eϸ����gmfo��=nt��Ob��8���9�7����B�P�E�O�o���ϲ�<�ʬxQ�����g����ދ��;�������BM�kG��6�ӛ.tY~��y��}z(W1��5L^[Ȓ.��]�K����u����=v�(��p��uͻ���P�t1�ZE�!������/Q�iR��L"AwGKwC�������^�����ۛPe���M��`#�H�fW�
i%�P�����@e���3�W��t<�c�ˠ�0++X�y�����6��!�Gw�|� �J��A$a���>�v��d� ��#,,JQp��^pW Ĭ�)�����POu�Q�(w�pbޮ�ПL&�Z�(�&�����x�I@�Q���/�#c2�r?+����%A�rF�R����w�?�Tg�r_�������{���=�_a�V��������o�`��~|���p�����0�CK
,�����훷?e�*�K�Xʝ��.��E��� B��
��|���fa��#M�y@0�	�K�Y���w A B?�T���v�F<�K�$6��=�@:@�	V��o%D�o|r�ѡC�e��vww1�E�iǓVj;<=���w<�` lQA4�i�� iR���2�kά�N�"ů	�ϧy�Q�')�]{��'r��{��/�o����8e}����,C��ׯ�}�x�ė^'�k ��O"s��Q!����?��p0�z�G̬�F�b�!��捛���(�}�Rĺ��E����>?��cb�xHP���4d1Z#Djӛ1�� ��� 
*d��i��h���ܖ��/Y��� Jd�Z�^�J_gy1�O�OC���75̌$�VO��tc]t{����1
�B �� �Nr������DS��|�9���ٰ*����/�����_��{�����R���ܛe������Je����anXB��V�L�.ݤ�}�k���/'�����"��&��K7�����^f���l�|RM/���>���d��;��t�kr"b�I����Ͻ��7����6��c�i��^��ۛ�9礎H �Ci��	���pN��+A�����o�e#+�z=(V �'�@!���H�5 Cf��
�DP�i����K�C�Z��i�_`��}�O;V�^�Β ^��|�p.@��Ĕ�<u���ܔXͲ^Rh���a�;�]"�)�*�7��?�I����[��9��~�s_:7����)�YGH`�� *]�w�p���?V�S����W���N)H�3I�TJ�g����>�v���x"��>u��g�(�>92Y��U���gG�Q�^.���P'����R�͓��0V�Ƙcjͽ�[�J��������8�<D<z�>|){�� �d�<�)q:<\<�`f���wr�@��QH��
|q�;�?��F>2sC�S�ӌ�A)���p/�[� J��×��>e��$��
1T���DT26:)4kd���V�@`o�W��2ɏ��k�Ի�V��W��g��P�������vP��4���f����C2 r/;?�hP��I����1Ed�[����={��IZxo�d2��Yi�t�w����;���GH����؟������"�{�h��*Vױ_�'+�W�ui-m-��b�r�#�p��<����&�1a��~~CSt�/���ʗ:%!"����D�Jڃ��o9sx7t�p4�s�C�Z��&�{�9�4i���q�� A< q�}�$ H�$9�Oi)5#�T��Q!��M+WlV���{�>��}��
�4*Y������ �2L}�x�2T*ػi�6�֥�W�+�[���p)B~2�j�?Q&aEdX�`�ɴ?����&��I����s��ō7�Ĵ+���y��\�?��m��3� �<����X����8{�,�y�\�y�|�<�r���w�܄1�Q�݈/����')�ە��+�< �k#8 ����Ȥ����СP�#�w/F �F�>��H_�^��\ 3��Q�0 �p��H�N���'ȳM�g:'��wΏ��=���Ɣ}3�� <�T�J��t���e@B�����Q�"�(HP�(S��?��2ڔ�ZUي�D�����Z0�MgG����V5+N��~��5vww!lmmaV��Y�&g�v.<���ڤ�6�z�hU� ������/��,��;��;�i�,�2%�u Gb�s6�<���!tu�g B�����D)�{�����Y���f�CT��t6���;�B �}�[�����5	}(���q��*O�.�N������Qณ���;<
����ó޷��]�J?h"{�`�Ƈo���so6����G���g�I��$q�ϒ�F'�}�[>���r���R��|�����}��خ3��ѼDf>-)?7�z����;�=��,Ͳ�F�C��J�� �B$"�
y�� � �uI����"D*(f��U@(��(&<	^i�"$��6+�B͊Ib�*#���H�Ib�!,���Դ* �\� �Z���Q��ڷ~���ج�1KD�̤�Zk=�I��,˰s�^���{�Lo�D����?�'��]���硲E���Rʧ�F��P���]���1�J A)�s�Cu�N��h��H�E�[աýx��?�XMY�:�P�^)�%L��"�A$�.H���A	)�B�7Q^�"@��h&�'��{OeY(�*��!��@/IRff�C<�V�v}�=��s�����G�^������ɓ��f���G:W��s�s�F��Ȳ30Z�9綈����.z����k��@�b��HN"���&�1������2���N��C���T�:tx���W׈}\+�t8�`"�s�9�e-.X[�;cHi�+�b�����;� >8�(xq"�A�V!��"B�YvΒ��O�S
���>h@3k��QJi���r�:�U4~xk�׽D���y>��%���eΜ�A�g�u�&�b�Clll�V��t�;w� �{���]�L�iVLo�?�?�ү�گ�����Y�)}�lr�f��mKfa�%�HH@�P���k���Z�[A��o]"���P/2z`�(m���Q�yo?f^R�����q�w���=���e�b D��B U��Xc�R��*Q"bD�/>HHB� A�D%�+k��W� +"�	�FR313)�t��e]�˺���b���K�}f/�Om����~���-dY���0�L����Z��
E�������o~3�~���Ʃ�-�������U���c]ҮÓ����Z��A�RXA'�����f���6�� "D�s�p|�:��p����C��6ډ��$ċ��z�ZnȐH�'B���\� 9 �&�q�ИN���i��b0��H O�!fM�}`kmduPꕣ-/ū
ߊbȂe�W�o��hI�ॗ����3��bVL���I�N��:�1
��֖ ��Q�=E�� p����_�tx���>}�;���Z� �L��D���L"� @���]T�����^Glj���*�{����ѣ�� �(����v���x����:Q��*}ǭۼ�>��<*�)��ޤM��"���dfx?.�:�13����i�I��:Q�;����V�ݼq�{�(�,� C�9sÍ>f��s��eQ!� �ij��A$yֻ�on������S������H�]f�ƀ��BbK ����zi���0F�V�4�6s,G_�:���Щ}:,���I�����!e-���z�!���2�h]Oo��kq.j�I[J�<�\�&� �M�D������S��E�/�p���}!,����^�G?�Q�>s����-����j_��V�$�h�&߶3��s�_��_�8^0<�;U���p`�@���wU�6D+�*Q��(Fb�# �߹���Б��G7�u�P����Y�t���f�ZYRט�ԫӴ�a����ץ4Rjq����Mۦe"��UU+h�s��]�~8�{0�ϑ�9^{�5|򓟄��,K�z=dY�;��6��eY �4y���*���a���W���~�N��/�������rG@v3���l2�['N�����c�q�rVS=�L�&AE��)�$���CQ�0f���:���YO���,���]m���y���GᨴG��[���A���<i�`y]*�G���qT��z><H�����쿣�J"�8�����p���W�պH�"V��8LZ�|�^�m>h�i�u��u�~�w��yy)�М|�Fa���������.�3`{{���'�$��[��N�:�O�=�d��O�������+ ��#|/��F��W_��ߟwtFw��ǟ��'gI����I�M�1���ꢬ��@�A���P�S�^�`�F��u�p0����A[�jGyv}�p� m�|9���"ǘ��1�ͺ1�<I�4�x<FQx問೟�,^}�"���
�~����p��M|���&�n���pk�Iʋ��w���_}�T��S�zU��׿n�^��Q��J���Y�5��ΖU1T�9I�*ɒ���&676�@��$�,�+��l���Y���?�>��C�Ԣ�9�A��p(��~{��6-��kCD�A��Df I4�"xo��p��ŋ���ckk!�z�y�<�#�{`����0�_*Q����n}�W�W���_������Lっw`���K(|;�^e�NΊY��e���I��Ι�8��^�\�qeY@)�T^p�r ]����z=��t<�ѣG�i��������|���w��1��qǿ�$�q�A���D��t�T��/MS�Ԧ����㻿����k���ad�<yŬBUY��E�߇��wG�����ɫ�;= �_����#�P�g�;5���'/��3+���~K��D�S���p!����>qr���Š߳��P��$�;�M'��"(X��=�*=ݓ�QX���t��}ʎ����3�(p�>k�O���,���I��У/�1�����>}�}������_��!��41M.�9�#��R��z��{8{�,>�����q���:����O�<	[9��3L�%��iT��wn��	�N��?���<Ҋtx���J� �dU��
W��/�$����_*f��^B�C�~n@Ӽ׳y��T�M^���B��#�S��v���Ӎ���G{�����yW��t�5�>(b�~���j���+}O����s�~��7/��(�,K�$	N�>�4Mq��&Ο?��/�ĉ �z=�GwB����: @�|�]��Z�����v��V��3�V� ���a*
C��>#���~os��^���Ui�W�$K|pN)�$���{���F��,ଅ��������ĕ��Mz�U��;��xԤ�Q�q��G���Z�8��o>z��1���?�wl?��w����~�m�z�u��A<Z366�8u�Μ9����x饳x饗����(ב��Z��ޞ�����1�ͤ��{U1����tK�u�궹z����f�u���KL��`�����])ڝ3"٪`�[;'w_��˷.����ڀQ�0����1��?�N���#��;��?G��q�5MSlnn⥗^��/�������`���[����{�5��)��@��ۓ$�RUe��J��i�X+����
� ��}�k��o���1�L&��A~{�u�����~p���������);33܉���IY$voJi�(�f���z!�JA��^����&��8�E&�A��񷸬�q�\wIBz�N���#\!����*���8��0��m�0_zx���܌"���:y�Į����L��`�.b2.���9ݻ��r���Ǆ�1--}��k�5eZ�?� (Z^��}|��,�g��Z���o;��#/�9�bu�����f[X^�`������i�X�+����o�w��ς����P�˺O�:�q��n���s����X)8���[*C<G\ybu\4�,�=��j~�����b�7k˥v_���a9G\���2O���i�a���v���	/ƈѦ3Dc�=�b�Z/�)��$3�97Oc�X2��p9��u�=�ݞ�_�� $	��:�X���`���^�Ͷ�9L�S����g�;}����!@��߁swo����;w��w���K�� r�����ކ���wn!�����7��ڿ����� }s�G>r#��>&����'v:�}��Ib�щ�TU���$Ku���ΓىS'�k�����[��;{�����H�(�.ԄB��-� GY�c�+ R$�x�ѫ�iy��ݣH�Q�����p��I;~_L��'�-�b����v��U�О��ui�#N8���`��UR����#��d0֩MW��&KXS����H-ױٳ��X�4����q�:Z�i�����'B�4�,��]�vߵ��>^麜���O�6��y������m]>��A$pRH͵��PUJ��9"Yr��2���r�:�T"�l6��I�W�r P���>\��Ƙf��v����kκ����H��X�Д�Y7c6���hD���oږ��c������6Z��<�Q�2'ζ�^݆59�~1fBX?�e�܂<���ً�ؼ|����곤��]��n�Y1��.q �e	�666���1�q��-h�������&v�<��    IDATv^�Ω���
�{cTU��~�����>�*XW"MS���e	�1�2���&|��݅s3����W�^�z�õ����a���i��+Z�[Je}R��U�4K�,K1&U�1��z`����o��y��M�g�z.���u�>�Y�b ���y �����	��t{�<G�"<���(�������Ԋr�S�:��������-�����:�����_|�o?�Wϵ��V")\/�	��}���M�"'���'����j�����
q�5�)�q���o�]�u���uM�޳�j�����:�6n+AD�(2qR�u���*Xk�$YCļ�ͲWq�6���eu�c��Q-�uH��9o[-��QJ�Z�(j�,�:���&6u,��F!���4M�k�[%=�ǵ���^��4MQ�%��+�r�R����W�U%�M���^%�]���.�s���?��mߧ�~���ƶ�Jg��C�����F���}�6nܸ�,�p��Yl�z�?^����Ac6��UƧ>�=x���B��_�1��0Q]g��G�L�(�+���c_�/_�r��O��>�?�]G�{��o��ܻ~H�4���$�����_����Y�J�P�4�3d���i�ʻ���$�~�����y�����G`�B A 0Dh!'��Ȃ�3/���C+u��v�x$ȡv��S�����C�C��=����X�.�0����ww�q�W a��|��U�\:��~���)_�:��z��X:_�	#�����C�˽�������^���������th��D��G�������3N��2ah����{�Z��������2��%"`�8vՌ�&>��B�{����@UUK�_]�UHD��)�2��<�6̲���&�J)h��Hk�L�~Q��n�+n/�r-Q��&�^:.֯m���5�Z����`�d
o�z�s���kױ����n�����S헠uc���^�V�G�g��g,@�[��v�m���R��~s�i�$�%�~��e���1�
a6��Zcju��*��H����}{��)�Α�H��Z����PFa4�C�ll `m���eU�t~oT��N�������]�rep�ʕ������w#�c��YQ|S��|Wk��^oP�keU��ͼcDBe+�����i��=,��2��
��1X1���� ��C�jӮ GġESp�[�:v��y|8�'���k>��$�i�A�r�vB��a�')�`���^<H����O�,�@,@ K@@ I�]���(���� �

Pj�vi�������b�W2(���Z,߽���O��������ʣ����Y#MR6p������= ͏����ܨ�/J���6ɉ ���.�H� W�Wz�\��=��:�*m���*��H��9vU��][�i��/~��#�J^Y��$�L��,��i���ܼ-V3/O�(��h�����KkmC�$iHO���~�~��,K8�`�bY�$I�r��G��LTۤ�.B�e�<�ֺ���~�'��J� Sm�����jz���{��������n�����)m�3�IDP�e���y�<�e��Z�5i�ĭ�OJ)�8qb��3^#�����%��_$���J)8琦9�,C0��*��N���� h4 �n�� ;;;�o��B��{{�U��V(K����7�����?�?_��?��3W~�J��u8K� \�tI�<��Zo���`#1C����D��%ȧ��,K%5�1������&�u{�w�ڻ��n��hei�� ��H�A��U�C˳������ e=6i��P���ں}�(���G�i��ïϭ��dd�\m��uXU����u��u��:����Y�t�գ���quP9��V��^�7��J�	��*Eј�V���sr��t��a�'�֪p��N	)��2�V���:ڪu��M��HE��d��H�VդU��n�6I0Ơ,KE��O,�lV�إi�,��~o��\�d��Z'�WPS{�KhaN���sB �f�z�}h��,g(�
֖71� B�N��sq~=�*$I�$� �9�RcR������) !Ծ�����'���5��ޣ,K��(����Hh�ב������8����'c�y���m����j�|-�tF"I�Rf���9�b&�K�d�'ܐ�<���a��Y[5��K�m�m���	���}3�"�t�5�3�e��aC򫪪I>���y���w���7Bo���g���y�&n߽��(`�T�w����A�o�������_)�\��[W��ӻ�@:��PIP���3��l03'M��։V��}�W���<K��r.��i/�43 e��8�v�;��w����=�2�I� F�F3/���Q�*�Q��ㄠ��2�}|������"�>�?�|G��z�<h.7�N�h>�������7��'���Ѫ?�:��J�ڦ��b�6�����b����?P����0����^����>�ܹ��h��H�&4͹ԲIk����fR^%�"�4S�
���U��6�j�'N��l����T��6o�rEu�MҢ�U�H6"��L&�m������ �nUU�iq0`8΃K����F4�NU�V�r(60�Bb2$��V��BeKx`]	g������E9�b�43�����3i8W�*\�`t
m����MK�`a�<u+�I�Um�$�_
˪� ��su ��<�/<�C��G�1޳Z�#P% ��h9� ��i���~T(��h������Z�,� |�͘Q+A@��*��j�Z���.�����X��A�1��<�c�Q?�����ss�n嶙����gM����m3'�u��֪��c��������t�ɴ�d2���&�Ҽ���mܹ�k+y�����`��~�O�/~��~nt�C�C���I_<�������O���W�~f�+x��!ȧ}e_~��A9����:�]A������}�=��aooB\��5~}��F���aJ�B��Z��P��}�v�O\�T�'O'=G�(��0�t?8�x}��YM����S�$�e��k�LŴ��iژ�bPF|��f���Gr����|I9l�mSO�H�	b��_"k��ŋ"��<jD����qRUJ��YS�U2֮�AJ�`�[�O������گM�������?˲l�Ik<gUU͟���`���~��O�UUa:�b:�6�9�&)'N�X2oF�e5�&��H6b����`{L���n�]����Idiִ�BiT�/>��Q��D��c6�-)�JŔ/u4�IL��&��s�9�9)��Y)ds����x	2'm����$s���n�f������Q�Fǀ�,��=�R & ���ʞֵK���KY���sEQ��k�8c@2�Q��8�G�@X(�޻:�̼O���b�<��4m^ʪ�p0��j��E��e�,�1>/b�͊1��:TU�J+mS���צ^ ��_Y���Y�������Y����ǰ��N�;ބ�B�����2��5��+��g����>D;tX��"} �˗/��D��>m�R�n��}��R�7�?jg�~���y���i��F�Ėnp����ƍ박ŭ�w0�`t
cR� �a��h�m��ќQ��'0F`��U��c<n�S)��1�ALC�����SќI�RY��H�=�B���n5o��r����f�iO�q"��/�!��=�k��o|�����b�g�T4�O��`6�5���(�E$8q�h�h�����v�^u$oO���%B�$	��>Ҵ�o�6FD�B���&�<�s�Q�vvv@D�lM,�/Sl��O$h��i�6�p8���.��h&���Փ4M�RUU=���7f��p�`L=���]���X�����4M�mj���� x���`&��cL������ʲ|~�rZ�����B��&�跴��ь���Y��r�ǣ���|E����Z~\2W^� �^��c���e�2�n�:[�c�/����{Hu=>!��=�E�F�Ў�m�x�R�y��o1��DP���CL�R���ǘH�3�&��eH�UY�:���<R�ZL�$&i귪�:��$�ι)�&����xi���\��u�������9�<���	��s�u>�P�~�ߐ0V�o���
A��?h},"��A "�����O�⠈-)� �>Q�E�v�(TUiʪ�B���AC�� @���QPJ��B�i�".�(��t[�V� ��%`�"h4�U &��V�����?��~.�O�. ���Ν�鷾�.��r��+��x:�_ �M<��}g����/�ߡ�x��/^��_�rz��;����`��OhCQn�E":����r���Z��t�1͒�x�U�0OQ��Y��x��N0�0)h�@`�5�Q���	 +��	L�!XW�*-�^V+���<$� ��P���i�7�j�@[-h+�A���1�����;$f��,�1?�z�F��>Ey�7�0^?��C�e9Z5q�	fkk�1_E�,��#�&����s��lS�?����S$s1:��NTVΕ�5�iH�s��%I�y^����	3*M1��s��h������M��bT��|T��m'�8�Gu=/�}!���X��9�D��M-�M������*g����TB���OE��&+����T�t�U4�IӶ렍��,ʲ�u��'��/�[�H{ۗ/��2˶�p��+�;�2�Ib�D�67�y�a�J^$V����aE��"��W.��]z���lU�HA)��F����0�`���#��|=�����C�j�"�B�9�����_<��������ypZ��jk����ֆAP�}]��Kkh�ʲ�1	B��y"q�	�X�֋��Ԗ'�� !	B�P���&ˊ"DD���@$�a9�IZ�Ê�3��z@>t�\����xϹ��x 4��$}+R�BX�E�,�$RJQ����2O K �CL��9��'�@`""�P�EH <�aR ���zAsP�,+vD��k�l! $̐���$��I��;@"A��B">!b�U�+b��Y��_��	#d��UT��t����ݟ��y>���?�L����A�  �/_N�a��]�PN��O���*����dF��aY���a�;߳�K�,�$�Nz�0��BH����N�X�QUD�(�i�<O6cR� B����ij�ۊ^�,��A�h�icTs�Z1\�����تI�p8�p8D�e9��"����⧔�x<�p8D����d2i�^���<:����l6����� ��d>��n^��R��ͣ����s��\�:|��R����a�##�"M3��1�ჯ#���H �4C�&K�l0)H��6�B�#&dUK�.��AԘ�j�!����è�(�k3�yZ�������o㱝#��j[��8��<k �s��E�uDg�Ӹ � ��R�pE�)��lND#q��D9��s�U��¼��m�w�?S��ڼ��^ӿ�����IUU��!oT�73; ,�T)^'�+�l�JIT�j�#�I���/�H2�@��+"��M~��פO� "�+�zH�E��9�HC)��0����yP�dA�h�l]pD��5�@��H�/����L�&B^���y�l!^+dV����}W@,
�"u�w�y�uU��^o���nN�4���LJD�H@�S� �'"$@��Je-��*[��2-�����	@��J��r�tU@��HB�E�D��G�1���H $�A�AAI @������2 ���sW,AẀx�V|W@=fQB<��D��$x�����)	 1	D��f"�~�pD` 3�ibė�kbH^)eCDLM�������(2b�)E�$�'&H1Dd"H�2�� U�{K�f���Ay	��#;�wn��N7�����L���G60��ߴ �ʕ+-/�>��7��{��{�0εҼٓ�U����T��,M�D�t��̺��?���;�ub��^� M�4�$�xv�Bو�H��677[*��RSTc�!�m,"jT�����Of�[2��sE�0�����H��&f����*���P�A��2J��%�|���H���KD�Ρ�*�������D�Jկ�<w쟓�:��CzC�S:4�~B��O$ޕH��A��{("�୅���5Rc�ZCs��! I3���ے$�u����{ddfݺ�MQFR�L����ؼ���K��z�٘���Jf$!U7Ш��k�����<����F�6���~9~��s����:�k,�U��)i	��{kG�UCeA0���9X� T�bɵ��&$3�8>�Ja%�2b�,_��^ � n�w�5в���-^�V�(�c�r �����Xs��3� ���{@+e:^gS��cV	���%�@�(ux�Zz���������ܘ���P[�}fh$����C��df$�0zD$]\\�܋��{I� `�,�ٶȔ��ڳz��<"Aw7���� ia�7my`�̨��XI���ԡ��Q3��Zދp�ʵ�#	�^m�������$ #@3/f�$�H��+uiXҸJb*I���c����X� 
@���5��v���2�e$�$4��w ʁ]2�sl�"C�Z)H������&�d$W	��=�Rmm	�F�E���g��$�@l�F	� pA}>��/ R�(���W�JZ�4��\�'$I�z-�nM�[�f)K'�p'�F2�S* D1 ����ک�m%xEr���&��##/(�'��mD��v&܂hi6��2q��%6 ��-�-V��kt2E��EDTAFh��b�w�j����=i+i"�vfv'��H�+�Y�h�����>��s���m������=�����������������O����T�e�9x�ʟn�G�/ß�c�'�0���l{r���N��R�����0_G}�a���uj鬐����k$2���� ��������G'���������]��a��~z��&6<H����<ߧ�: 뚫u] �#=߽��>������S�=J�?�ൃ�^ŷ�4Tv���NN6�˕�7N2�`�۲f�^(�nΖ�S	'n��ܐh	��B
�XriZ�h�i�D�� ��2-
����ѐD�	�U)�Ī�(Kw�4YA��&W��2B-!+0�2E��.3�����s F�$��2	�18��~��Ps:�fT�L��*�#�be)d��0���`BA�a����v���PI�̤����T�

4)�L��f㍹M]H�$P�)d��L/t/���%Pf�D���%�$#��,�~��\�2QA�R�^��(QS�H+���֖u2c�֧��@�P���}D��RH �G�	�_� 
JI��!#���:=Y n���}�v���Ğ�
��d鳼1"rE`�TI�)�h-/I��l�@b�
Ҁ0�М3cf���A ��2@ �4���3��h��o3�k*�F�SP����#���f��I�+tC/���u����+�@fJ���L)�H���QIb�q$A;%WAň!%8�;A'�m��  ��J��_)�KȾU�^���NED�7	�X�k +�'�8�l����=I'���6�k
��4'�Hy �m"�A��ɜ� ��p-��M�yVk��T#���nU �������ni �B��|&F�% M�`Or��IR��%��?북_��~�ܜ��'O������8��c�>���իW�����G���N�yi�+���"�|���T��t7e�Z�l�O`�֩�@�2ġ����x9�O���qdɎ�s>AB�p�Bz�f"p�jzT��ʠݛ�>�a���M��B�h�;�6��8s�������t�?4�P�5��.�D���H+�Yk)���$��Q��3�\���H){>O�{�ہ�."=�v �Q��)$�v�9�6�	 ��F�aZ铨g��Y�3����0M�v�XB2t�8����L;��׵���Ief�gt�X)����������}vP3�sg�jdP�Q�%47[����1�B]�Y{>-S�'�  �IDATϻ� �2R�y��Պ���80:<|�gEĆ]`�#���fB�}R �IY�$.��P ��́��X[�� 2W�Q	,��8Q$Ԛ��_�֚�e���fՌ�nT��[�sR�ݥԤ8egD 1��"A�1��,)A������3,(JU�$o�>$��=2�Hj{�5�M����Ho� �a��!�*�$�9�	��-�;�/��OI�SZ	��䒉;%�ILNlEn��H�S3���]n3󝄕�		�TK�#һ)H6�n���Dx���^]j��!͈�Ɔ�J�(ak�H����"?��-3�B�h Q%��ߴ��ɖ�7� �L���r�\�]�E�B�Uٞtɥ"3P%x,�=��@��V⍓�('U��q�d�RH����+��{����Lc"E��\͆�\���U�G08����6Rq5�F�3$�L�-�&���*�+w4)���IM��t�w�ߺ#����$2�-���5�朴pG��(�� k-�k�gt�TgH3����Ӭq���f���&NOO�f�������_��o��W�^�v;��x���g}@�Ꝧi�L_���6?����/�C/+��n����M@������8��$Ǻ)uܞ�T��m;h,�����=�8�����ﰎ���x��#�Ɍ#���*/�;�΁G �R��(�`5ph;#C���PD�A-"��A�:�$W7��-��Ks�=���*)�fls�w��T�c囓M`-^n���m$�������m�k��[@��F"�|]��B2(�P�d��3�b�������ڕEY�|�wo�͙���s��O?W�g@:�4Zs�5�W������L܁E�H- �N��WI)E�Ҋ�eY���.J�p۠���!` 8+u����	��n [6�͔�kk�����( ���x5)��x#q6b�Y"e,�˺�wo���,<!yzD����~�����ȑ�9����ImP�+	; ��!'�čB3L����aߦ�Nfb/a!1H�i�:�`�"�k�)�f0/��~��Z���'f��r�S�l0�Q��s O��g����T~f�gF�0�.�k�R�\��݀�!ٔZ�^Hy��i����e���� .����f5	�������ߍ�˔�ؙ1$EH�D
L-���vR����H��B�!�s	{$/�!I5�A�.�?P h�0K��( '$nIJ�(J$�0H��n�_"4���쓐S�D�<S�U�Ud �A@��um��+���\H*"7f~����R*;;�R�LH�6������d�_|�/hȬh�$Z��R0�h ,��KDld\���v�kF��b�j�Q�eb|)Е���
V4d{Lyr�zY���� r���8��` �%w�1ǛKRb���ZaZ��5
IX+���4�P_Yï2��L{W+�Rָ����zJ��lssz���;ȯ��*�����=�w�ޭ_}����k�믾�˯��C_8]�����_���o�����������_�ի�����-��|����EU��,��Z��0�i�4����8�G�mj����A�r"Pͬ���D�ѕ �g���, ~H�t	��;i($�~�F��9�\�eCGx7� �M�i.���  G%52Iq��ݲ\oo�-3��:b�1��p�S�F#�&��*����\�y/7F�N����IO133it4�\D���)!�{�M 2%3���fZ�"��г��֊�p�EȚ絖��g���\� ;�� ��s#��0���?���[Y��; 3L���\��d��-:��.h�0)���7����D~"� `�]�R#�~a��M�|
�3 ��ncm����	����w�~���1��k�3|������ߓ� ��ไ3
��wmk��.)�q߱%�g����i��c^�<!��]&tA����[C���F��F�fƧ��<Д���_�"��(��� |�@�X  �[%6N�*�6�.�$h� �=]��,�3 �J���[#/	m�)��4�)��ĵ�Sx�^{P%�;�{�F	���m�.�ې(i�-0p� �� }���L��4dg^nL����܆�"�&����r͑կ�r�(&��y��%�;I7�o�	if����\R��D3�-+�%z� '@[4��#y��}E�ȬP���wsY��G�Ӣz��f.w�����Z Jq钭A`�{� @�=؈@9� 9e� d:k�{[@k!��� �sRՒ3
��C��Y���-�e:��<���V�/(xZ��F,c�=��Xչ�7f*)T�eڍ��L|6���ʥ*��lD�(k��������>�Э����͛�>xSk\����Zk��� �Ln�Z��,w���`!� �Oc�ئi����NNv����z��J��>׻��ś/�͗��իW�c�������} �ӟ�����nj�'������l*�_M�|�����?+�gn^H�����͆�1���Jq7�.����5���I��3�� ��@�vR��� *�VX%5��A��4)�̱��W;�+׌Ʉz֘G/+	2�F�5���ܴ�g��ˌ8����R:3c�|ۢ���)�Y�&h t�n�ì������V�$9�B��.�fU�W7��Z��P�@��:��eYwkks��9i3�k���^~'e4(�	��כ�Dg$�م�B�R�m��	If�
�Kwvyf�8%���N`lۥtr�� �EK�]223�Pb��zrL2���R˥�C�ŀ�T.���v��D~"�ԀJC�~)7�)u�J��h��%]��IFP��Ab�sr�����$]>��� 3䚀���� ��Ժ��^�|U�%8#1��B��̼7)�N���a�zuHK�c�dy�	��.�*��	W����Z �t�@k0yxfJit }�?�?l��g 0v�%ݍRKX~fBK��akB�H	)�M��Q�Z��_����B܃��F�P&ҽ�݅�ѫ�#Jos���M��R6���um�R�ko+9M�L�<��@����k}��w�����e�p��_ʬRF��MS���� ��d���q�I�vw�ֺnطO��|�u��~��N����z2 �ݨ�:�o?��D%BelH�-����C������,�M �>��0WL��^�]U���YK���sؕ��~�eZƉ�ɾ�����%�' �a��4ޞ�v����[�8��
 �6��n�?�=����˟<�����ܞ�ɓg�!߼�B_~��^��J/_~�������c<�s�AAЭ\���FI�M��fu�/	~2��8����?+4V>#����W��҉f�&���TƗƣP;$n(�ӱ5b��LI����7�HQ`V/�(R *�eu��g����dH�h&5>K��id��t�����
3��NK	��B�����
p��0W�S�߈�4�M�U H����m�� \�-�u���J����q;όZ��kD\R�IF�>y��-���Z!5��D*$:��)0� @E�3�mf�+RA���$M�}s[{i%uH�5E&��x� 3����DO�Q�" `�`�,�0�JQf�J���
q%R;�H{ �������$��0��0i&	���̔��y�����L�d�(�/#��.����.-���(�@���i��?����Z���³�x�̜N׃֨�r`g#��l�ZoKQ!}<XY`YZ��eo-�����E���a ��{���,�e9M0��Y}y�o;��'����uX+[��� \�8p]g�:>Lo0σ��;��p]��6��eYUʠy^u�G뺰��q\8ϫ��է�O�5 ,֥!.�fX�}[�ۍ?8��k?����у��:}��|�߾̇��>^qh��ǫu�a�t{ sð�_�,���3w�u/,}�����q\�����_���z��<m�������.���۫~-oa�ߟf٬3�s��f�A�����(Ĳm������ v��w��x��W?xN/_~}��ի���6� �1��?8��W�����o���nv�� `:�k��,���3񒴉�k�Of�A�_�`@R֋1��=L/�Lu��ƍQ/H���{�P�&�)�\�͸d�dC��� �������U�p?�Y$VB�LUR��AO?1�i�ש|����h��{ !r0 �v�c���4ebDv�����(����1���=]�v��,LLh�AQ$Y�7�|XVZ63Xʰ����_m�h����|5++�A�d>e�T�<3��ߊ+���d+��%�V@rgƝ�-i��ꆖ�Fz�֙(��,ꂺ"�6�`fm�0��j�)V_�դ��=f#
V���'w�hfvkV@������fV#su	�Ze�ȭ�uW�����꺟5�Z�=�N#����6�~Ts�Ojp�c2�NO�ED��:�v�SEo�>׋����o���>\w\���;}��x��+�˗_�͛/���� 8nw\����a�����_����V p~��wi���i����xr�A�<�	<�8���7�{NS_/1�a���S��ސ��Jv��ZƱ��c�����wG 8Y>�P�f�q7�=:�o�z`7��$�ۉ�2r��sYfN��;��$���fk��i��z���V纹)yz����������|�m?γgo���}�;��O?}��	h~�K���ׁ��?�^�ze���ן�>��9�����5��_�����_���Y���>���1�)����c��V��4�7c7>}��_��!�3酴�3.���XO�� %�ޘC0 TB'�vNh��7���[*�tG�^����L��>�N�>�&F��pD&�P���mY��g���,׶<s��B�+ɯK��� ��xY����\�J#'4ݑXH�\[�@�j�[3�0r=T�Z�Յ�ȴ-����P�����9�8	��3|=d��^�e���ζ�"���
��b��a��E���R�KQ)m�`�9Pb]�܋�|�2oUc�[����<�P�ڙ��� �8�pW
��K,�iXі�2�h��ke����9�$����\d5n�Ǫ�o�Lӓ��g�a��cĊ���E;?ǰߣ��5����\Ob�R�6Sm�5y9_\<���Rʙٮ����N?\��!�t O_�9�ޯ?=,��^
���k�3#o�>���#�:h�7o�����_~������a[�3'�u��x/_~͇�>\��s=�{m��7��9�`��/�!^~�/.��˗_��GV���ա/� �1��4����O^ճ�����~:n��$_��!����2]��O;��Mf�@�!qE`1+����^�]| �J����N�v�׊�V�j�½�k�rH��)��c.<JA�>V3���<�}�2r&=��x+"[]��W��*��e.�e�(�ԝ�<_m�mm�4�-��,eЪv>Ȃ6S��tW�ڗEcC)�J'�9xk�9֕��4u��a�0�˲�f�����Z���C��I�]����q�����,�L;%�%�\{?����9PV2^�Xݹ������n��2&�I �d���6��%6��X�^e�s4�~�+e_���f����,���F������v�Dggo��_�;�����<����}��>\��I���#�x��x��x��o���> ҽ[��ۡ0W/n���h+[8�+q��iC��Zc�CT.�ʗ���G�0���B����S>%=2s��P�P<5(s�b��t�iLN�g��+�Ĝ�����Z�s[�7m��c�
 eַ1�S�=���|�7�� ���0����nW[[��C�J���t_jD��Ϙ�%:��o ���M��#�u7jwW�r��"�g�%�m��ۃ��+Ǯ!��>��`��lnm���!��A� gg�����_�`��__�_�I����<���x��x����s�Q��C�?�i��ؖir��l��"���Ɓe�lM��>�q��u�6 �����ף 9[���ib���RV�y��\� ��]�W��Y�Png-ۑ�Ǝ1�4H��q�C��~ G��t���@tqq����_<�A�c ��{�ꌞ=����~��y�+ �?}���<Ԁ�P|���ݴ>���1�1�1�̠�a�'?��}��%?}�������/~L|~�����ы.>{�#ktd��/���x�� �~&����~3XzD�����������B��K��    IEND�B`�PK   �x�V��!�D�  Ԟ  /   images/cf2dd1a8-295d-437f-92b8-7fcc138ae9be.png4�uTT]Ň��z�iF���n���n���)���fH���|k�e��̜{������މRQ��zM�a��J�?c��4�<u��Ar�b^�+]޹��<�B{�������\�K�B�EБZQq��SH�y����87�����o����b_�,��9X]�'�O!_�YM�cMO�S�ր���nS�[#~'���SB{��7���	"ݚ�g��)L ŪU4y�����[h! d޽�v�YHl��T|�S�F�>,��	�Qr�4Y�@>�T`Kc򆓓3�����=<�$$$�?�dff�°Ȧm�A�\W4�^l��r��!S%u��m�=�-Uv�q���)$%�_k8���恢�u�����G�j!��A�(g��r/���n���OOO��\�H�ژW��}���!�A���b�ԟ�! �0�,~*<V�i$o���=_���YD!�rL�ӶyV6�y�Q��>�K;�MV�+v�3�0-���c'1�] %x��8��������.F�6N�6�j����N����L��z���D�u�����ဂ�Kh�#�R������۴Ϝ����Q�J�w5�'�TB�G�琄����q��|����ٞ\9�s�\Ԟ���A�AEA��s ��Z5���͟���<s�P��I�̋�ƥT3�Xq���fFZ��d�F�h錓��Y]����A��ur�bR�n�쐝(�0X<(a#���Ό��Zg30�2dq���ai֭��N�\B�p��n���M�ɴj��$"Tޥs@�a}���(�B�3�����@T䘘����gs�@?J+�&�4��@~a.��au��E6���"�s���s���-���u�n���b�g3d����L@z���L�͑�숀r�{��͇5ua��p�����52�)���~I�ό��N�x~,����TI$qɁm���>��,�4��_:��8Ej,�nT,�"�dr�3���zmj��(>�>5Z�7�}KK��,��y��U}�8�d�ݝC	?�3U�9�O��}&��̬,1�n4J�Ŧ 
`	uk���%��#Ȟg�� q3�(Q��> -q�:���Gq���9����A`��QG,.I&���Y��I@b�����]鶟W~^
��a�����O�	�镏�~��2Ţ��;��������/}���;\���-8f��v���0���������U�4�;d�U���h�OK����L�/݈_��)N�"�'��!N��sFr���i)�i9���I@�@���5�8�ۈ�|*;	ѝ`0M*hڂ�PNX������M�Is���N�����a}�������ڞ�(�����`�5���X��هl|��2v���N�feC
R靾,�X�d���b�J�>A``�����Q�F��=)f5�������kd�3?*|c�3��!��(d�(d���Y�"c��2�����W3N�+�Ӻ��􆇯�)WZ2��حwSt�n�`��
��u�&)W�a5/�#�� �xз���۴ח�_!��y�g)�n�������GC�I��qԨy?�ZS�WB�R�ꝓ$�{!X�.��:F�!nn��Pξ�Gbl$V��+����N}��N}_�P_��Ȩ66{�ZO6�W���J�GMmm_�I#��ˤ,UJ�W/b�I�YRx��~UG�u_�6���,�wan�ɔ�2jŢC��D(O���;]$!���Or3��.u9�./���=�[��u�^'-�6T��D�?�x~��H�/;;j���5�R,M��ݵ/�	2����"7�掆�G�M��}gI�j���1m�l������m�#����|��K S��JJ����tV�fqZ��f��<{�x�{�o�D.%k��76�Ag�LD1_Y0�ˋ�j�eP�8GCVqY�0�!�o��o��9��d(����YU�s]�tY�~üxB+o��U'~(<}8��zN�\�a���1
�ơ\l�_���4��N0�Z��p_-Y��Oe�m�/}��2L��6e�N������}7�|�v1�m&խC��|0��EI>�"�j�6u3�B�[��p��� ��F�G��AB��w80@�^K��;�Z�g�K��_n�$ɾ�qӭ��1i���������$HL։�� �#�,2F�F�	$�8CB@���ʧ*�q���G{j2L�UZ'A�����ۏ��=��m���Ï
�o�>�XB�����q��k��K�h��e�`�aэ�ܲ�3�` =�� �"��օ��������T�lwq��T�l�,.��h��樻,�?>�?Q1���Ԙ J�bvjD���i	�$�������Ӓy[�4y9��Ye�����
����nad���;o�(80qF��� :�c�ǁ�YN"7�ƣ���o*�ߚ��"EyQ07�=�Gb͏�dc�g�3��gB'�LJ�K������W���͚�46
&��H�Dwp�}���R��{+<����,9������݆W?>��p	�š\4BH�C�83�#�\�a(fP�8t')O�3Fn�t�����n�H;.|�uE�P*ư�v�Wn#CV}�PoΩ�	Ҫ7dm ?��"��4����yV��ʊ�$UH��S*j�lWM?Դ�l�V.���]]]�yyR�I�%3@T��<�P3��c2z�BN>8:*{%�{��8������YU���N�twƞ�u��9j�c�{�t��B�ȑ-\J�1�60��7Ev�O�rgreS�$ޤ�I�"�����SZI���B�U-�ۚW?�ʱk��l��lD_po�� ʹ�q�ܔ�~�J�NCo��8��!x�Z�,Ftϧ��̜��h�w`M�������"�uT��ONmB�����gm�Qx���L�c'�\>����Qt�7�[�\�MH6V^��Y0Cq
���a�/���F�4a���B��6�jX�پWTV��\��4Z/\���p�*�r���sѬ�$�u2>��9_D�mp�M	��P���hgc��QS�u�kӍU�;�
ի)Ra�d��ۮ^8�n����7�b�L
�jL�N��x�Q��{����5��*�>��M�����oEҠ�i�T�%#&V~�T�ږ$O�m��H,��`�z��;ޙ$=�~x��g+���ill4�-2�Wx+���ǲE��~�#m��co�E,���T�jo�v�xa�#WWW�E��;��yX���ԝD��Xo�Ir[w�ղy�g�V-Kjڶ�:�܂�Yy*c�9�T���	G�����gFI��B��+";�I���ݳ����u�I���������|Y����(�ꆎ�Xl��c�gvU����v�90�~�V��5�X]��)f� ����l����pP����rwK�U�,x�J�}Tse)N\�2L�n��7�m�&�z5ZE@6 b �dc:�/d%u��C�,���f �$'s�<O��-x>??�Ƞz1J��"q�L�/
���r�Vl�X�E�zÐ�3����@�1��e�H׶C�
�R�G����]���z��$��rgٱ�n����I��^"���,B������~�R��x�rʲ�'����.���Ѝ�#+����՞,K�A����G
��pԪX�aE����4�mH�w�o�Wݴ"~x�s��Y�Խ3Q�[[�Ve��G2��-^L	��C�i��Th��<ʜ�zl�_��B�[�+�A�������}�i�$���
d�� ���>l>���$��)muj0�lG�������i\
�������%��.�]N�c0��	��S�-(���"������hHj�i�4s��8}Sb�<���R{I�%�&66m�8!Y��������MoJ��a��Y����X�覤�X��n�Cpmu���r�m�]B��=�}.�$�U��!502 a�Z5�R�uf@�L��0*�F�q�����[�$bmqm׬`���ǳlrّWTR�sb&u�,0߀�C�C
�q���}���(��y�G���[حu�X�{3P�qzS��8�O��&$ܰ�Rb��ȗ�p`r��Dȗ!��O�{�#�?[ф��l�ޣ0�s���z:#m����*e��pl�����)ӥ����'f�|BT>�e�7�a}��w�}������ԉ���*�;��N��R rOU7���X�Z�,-�6z����2ބ�-,���̫�jq���7�iR��֦7�����_�D���[3���6���!�73�P02�������|}�u
�!v��c�[1��E����?{2ϻ3S��w~�@�f�8g��*[p
~�?���	�:g�n=����)���xj��,�p� ;�ɳ�����_����MS � -Kq�=7��Ѩ�߫y��vk�
)bl��u��y�����Yh���WL�5]��%"Tp-��7�z���,�m��W��^^�_�	N�PS�*4���U��X��m�FG�95�Ь�̐2�	/
��.0�vZ`le�-�I���y��p\Qυ�2&��0tt�1#1��i�C�(�/��ю�W���J���F�>�"�4�_��L��T����i�f#w�&��ۨ�$[ɪe�;�W�(Skӗ{QP�2�S�?ł��X�]bz�Dn��;�,�L1�~0+��h0��F�/�k��qw�,摫�Jj������P��*���o]F�2�V7ց>3_Nௗ�N��"��g()�*\�>��J�SG0���H�v!I�Eg;�I>DQ�bn�Ji��!Ku���Y�d������j���D�s�@�̡��~Ϝ�/ԭ���B��>��~��U$|�r� f��G6��`����_Z�%9�ے��Z54o�Lc��,��8F����@�ov�kڍ���}�n�7bV�]ˈ��u�I�$�_V.��*�B����/�3��aL�,�c�g�y�[��^U�?��ـ���t����6b�C~Rb\L 2���
��`zc��~p�A>�V��C��W�}1:,M��V���y�=H���B',�Qm&�V�{qWCB9�T�Y3D0����ӈ��ٖ�,�:���S9�hW�J��`�P����;�T�}��6�3<��"���,�s��X����j�*Q$E���6�(�#m��3�f�.>ॅV�>x]�z��>UT�6�c�C��Q�錉"ެ�]�I�CCLVF��"������l|$���C�_W�?dj�.<��t-�:j�g��qde���;�
�ߑRŅ
�h�T 㸓C��ڸ��>�]N5l�S��d�����˲��D�٨[��?H�h�_>���V*H��h��u��p�u9��ˇ:��fT�E����Qh�^�/v���0�H��1��=R&��h̦¨�0���ƿ�0$�/�*�)QUj�}���ivZ$gި�	/��0G9{��3�Ӎ�@�T�Ҕ�������H�F�|g� \��-�kA=xl�kh�<�],�C��6\$O�n��j���!�U� :Z� Nx���ǜ~�Q��^�4GiAJ��h�<��`$����34d��-l@�6~U�+�|�b��Η�7��/s��3�,��;=e��\��@ 0��;���H�8dRh
.��ؚ5�6�Vr�D<�n&E�%OR0E|��o��y(�q�~��d���B�xm��[�,ܤ܎CB"Ȍ��==�����gDo
�"��q��]VqrX�֎y�����Fr�?ڒb�>�[�\��*���WK�~H�Ҙ������^�{�K��px�	��V�5�
�W	CN�YVb���t=S�Ϯ�i�1���F/>�[���	��f/Oh�r��ʈ�������i��oQ�;�x���yi���o��f���L�ypှ�ǊS���[��T���u8���fAp:�����I?vTj5�V���~�T0xM����{�I6TE�me���0v�z#g�I�ʟO�GȻ�R9�Ҭ��Q�Ar��Kť-wF[@��6Q �#CQ�s�"A�a園�ȅ63�z�(�S�u� ��h������7���x#����f�,� p�Ug���7�J+L��TGD7�b˟���N14� �����:�\BQ7���C2��C��c~�����ɯ�V�Z�>�g�X	��A��4J�Am۷����Q���/���A�gӶ �a�On>�A��8������ny�WhT��w8%����IC��D��0�	<��tt�`�<�.���/\WoF���|y̭��t�d��V��]���w!O#<�o�]
4�Iuί��oP&@��l��[|U�=�C�*�z^;�Kժ� �H"m[��l����5����M�o>݇����_��� ����P��c/������Gk�0re&�+?��4�` �զǮ�+��0�ơ������[�Pl�oR�b��i��Y�Z,����Zy��tqE�F2�tvâ ���R!3�@�5^{Vt�4D��^�̭̇s�����6����W�6�k����]c��A��q'F�>��-�K�ul�F��?��C���v�R�J�ίVE�U����Y�/��s�����$@,N����`�O����Ԩ��uG췖Q;�#�SңM
������&��fK��V�=��u���`&;����/��~zSV=%ʊ�=���'E~;���͚(�e��b��~���ћ<�<��Ej����йj�c۲��ݡ/;�g`�����6��ӧ�i�h
�<^pe���$!7�`�ē'��\[3�4����5ۦ�7������[�k]gIL���l��K�v͂O�C#���!^�BN��pAB��s.���ky��y�Jf��������.Eƍ�%'�m�$���7f�}7��^�w((>O>�-�!��Wa�L6"�(���f����%i�D�$W���K��Č�z��L礊�КW�Eˣz��x�P�\%���·}᭝�8%L����~L�6����u�{=�XE���NiႏJJJ; ���7��'�����-d��x�����?��۝K�����]{>TP=oܤ��Qx����q��a�<���|[��?�ӵ��?b93Zx��T�I]��b���뺊�oaL���#2�q�E�ޅP���Ý6-26o�bF
�}�:/&C��\}Uz��3n�P܄�7)�Zt�u�e���Ĩ��]Hw�P��r�����;N'm{�g�2�/�k�Z����L�(<O��(�8�׎�mOX˭���ej3j��]��:r�.������?82X0�^Q��د%���Q+����G���x����c������탊CכUO��Ӯ�gU _i��WV>�F��l��N#V��#�W#��3��X��y*�U�KWi�7�JX����V.��\�j�bj�I��ˑww�PR,���
 ��o�|�w���\�\�E���x#F��q����<g͕��;X�`uQ��^��T��������g�C���nTO3TO��-L7�K߆^q�u����k�����z�G�n???�Ӎ^u::��aн��g�	ɎN^t�>�k�a�҂���'���U����cS#%" ٥/��*�$x�/���2�T=�۪:҉�����L�����zv,؇��:�nV����_�c�����atA�YKF2�4^l���!xN����RK�� ��V��gHA���Z��)�9�^� w�1�\�ы��[;:b�8TTV6��!���*'��eu=��h��ei�?=�1�8�K�������s&���AY�҂���F�N�� �����k_�K�]���˭�{޲�L��c¡�=��	Dzy��b̖-#�RJ0�j��z�:L՚���]:�Z��>�8����0�~�ˍZAp���kIL��D��j4������9V~��/��NWEEE��t���ԩ)ڴ�h��Ԉt�+~�=9y�ofVV��/�a�$��pIf�)�	KNA�ؽ�@�֧��u�����#~�^obC�s����U~���2O:���f�����W����w������[�˭"S{;�'��z2K\�I�z�u�ф�p��I7Fmn�x���_�U��~(����ϕ��*��U;�*�B'��i�i�E�K˱5~�ZD ��(��?�U%W�T��_������d ��gj�P�!N�D0
��&���`!|Qͯ��a���
�k7��'�"�1��!H�2��殓c0��>Iv�]��+Č]Xk]*��ciɇ��h�  0�g~�� ����J���{E�lf@�4�"���� I��4Y��=�V�F}������>5�Р=F��k�P���	Qj�ZC����� u�m:�����4��������˔&�D�q�s����G�{];	,�q��:����Q��C�Z�s��狗�&����h����CF�+���xO�l'��;MN�l��jq��<�W�!��H�Kf��ݥZ&���0qpƧ���S����a�m�;?J :��n9�p!���dj���/K7.�**O�����"F^���%95%�>�ET�t�.|@��v0���F;\�w��P"��tn�v���"Ly���s���.��%���^r�伐D;���5j.~�9���Ͻ�~�j�Ȗ�e��J� ��J�e\D*&��Q�d��-�c�о��B�� ZQ�K�I���
�4�e)�466=����
���� �+��Eժ7�1m����8��j���Pt�= ��>�`�r��e�bgʵ�kO�9�|�_�T+��&D�͟��Ω�[p�W�E,�<�K�37W��8��)ˑ�L#���lK��7�-��h���_�~~��GIôU�L�e�:�>��b��E���6@��=^�dN{]�0��O)?��'��c?�Н ��Iy}��� Иf�D��ԉCDE�7����
%pv��P]�/�X�4=^���?���K���4,�����]2T������TH�y5~���F��B��Ae�O��w+åMX��/���"48�$�E���*V|�F�'#̮Z&z������i�Q�\o5��<(x���.[{�2#��;kb� ��������!�~w��.� ##����>��%
����o)�Aw��)sx�_BL�edZp���>X�K�Z�a�Ί��G��F*))�n0}�f0�#S���fp)����^^��g^���O�?���>����_�7у�dʝ�Gqu���B��G����c�P��d>䄃ůt��Z��)*��n7#�Շ���Ǉ^L�P��/� �k���p3u�3�eK��%T���P&��ju���"�n"}��Z��J�m�IwxG�?����`�jܸ�-���pՀH0�2o�Y J�+ꏟ�S7�����U��ߥ��2}pX����Ϳg�D�N�og�t��3-�0�&�
��7��՚�&<Q������b7���E��>>�/C�	 "Q�	0A� ���������>n���y��v�s�*��QX�\��c�3��w�H6Ġa�병���=�I�����S��@_�<�|�a��D�(_f�I:�!�&���*�d(���ʞ�e���fA� �&��|��Ȳ~������a��/�% ��?>~�[��h�Ώ�Q�FYz<���F1H�؅���������9˥s�9њ>�w���8Z�Y��ϔ��i�(Z7�y�˔1>�w!#�ϛښYFyZ2��� ɔq��}^�8�JR�J�j�u�˺�d5����2]pNc��A�0�����5���>���~q�|�Z�DlJ��͛����\��_M>y�v�x�|e��-5Q��F�wA 8e���F��d��r�?�0[�3 �7/7w��s�Ոs/_�쇜�Cv��Y(b��L�}�l�+H��?F��l��G<�!��ɔ����!����N�.U�xΫ?"ՠ=�W�u9�Z���G�n:y���J�Mf���+��R�"J���(k|�|�Ǎ`$�[���ܴ&���P��sr��5�̽�����6�-q������X˾w������.��:��<TW��r���/w
��}�c9�跩�?�=�4kT/[C�:-N9�Mb�^�:����NS=�̦r2�8�ߴ<\&�a]�~+3?��;.��յp���l�ۨ��G+//'�p�n��U�DG�ǡ�fl?��
 2@t;<�/O?���ގ��/�]/�~�^<��+�*no�=��X���:�ẵ(J1�r�}�-�H<�?₷��WC�ڤ�\ ��ۘ9@.��			ٯ��M��((�s��t�����(sd������ʴ��}�E?� �W[gl7G/��qD���i�f;?Ty�P=V`�PL,,S[�(sD���}�Jo<���$ߞd�a���!�_󾢒��[�+�p'�*|(���ů6��랯�8��y�O����V�6�g����zo��aK�pU�;Ez<@��^FB�^X�������T�u �����~�W��_��R��L�i����L'��'�"����8���It-���$����\^_�Q.m�0&�:�ڢ��l6�w�LoNV�fs��"p����	�y?��|��t>�tDĵy#�� TTF�C�~�=.�X�I������d��k����3 �;�����k��̾�0�y�ҧ��7�ԗ� ������/�;��r�F�Ɂ�f<E=�C<NV��>���[?��AH��ܦ��_T#Yb���q@]	#gq���OC���0�Mg0}.���a����h�L�M�j�]�0�K7g�o��h����;���r�tI���z��[α��q�&�X��2���7���rs�yZ������(����d^���m<��e�V������c4k41��!\o�1c�W�j�m"G��0�g�7��Չ6�9\�m��-��M��Ι��q��Wˁ�4E��hd�	Sa4h|盝��J�a���|�JJ}5?l��5u�����IN�`H�����v���g��1�}l�>g�/�R�K�$V��<���,�VVE���`����ó��G� �O���N�?�N���� �)%�U�m�\�dϟ���q��N�ct����.ׇ��1)py<��l}���ە9��F(����� ���tx/�G]�謍�(V7r��Ϧ��q�u�|͎�{gs��&K�?�1"+�d-}M�f� ��I���J���Z6&}r��y���;Uzϑn�h �����Z��1fc�� t��&!��F�R5FF���9r���H �K$���E�KZ�By=�m>A�[_�MWf#���4�`�����ZZ�-�!�rDZ�᠋���_��n��O,�w�#Fi���Y�G~FٸG�Z��Α�U{�*QW��s����|��0!u|:���9k�O�λ�k>;�8H���C��"���X�ɠr���@��G��UF��H�w�<~����-�{ ?�A�ժ�|�������BD��Ԁ��&��~���G%w�dɮ����tM�^1B�jmz���}�"C���B4^�\KyLIU�$b�͏-Y��?n��DP� �$b�ڢ?���V}�G�"�0Ԙ��i�5�l%-H[y�\�l�+�_/�~q�8nf����;�;"[󳰷������ǂ�+�7���O��S��X EJ7hz�<������	�y��tx�*S�" �*�����|�����N����#��m����a�߆ B�9M�{]�O��s��Ȱ1@�y)�k'�s`� �"ʎ"�9@�R `�h9Ef)��h4�5󶀚qui������0����7'C���l�7/�.%8
w�AV0�>���� {F5�Me�`^���q�$n^��_$3w��^_�|���ֽ�V{0h:��k��׆� G��ȿD�/�]��?���n|'##s��rS ��Un_BG'3���٢�ע���ӻu څ>���ހ�C�fcL` T��L?��ձ�Eő֖ cU���IL��4��m��T	�����4�&��� �VΥ'�����!�R�a�����7���FY�g�7nI��s��ŭu�:��s�Y�,���}�'.4��Q�v4ub��<�`��1�dT;QP-�a�{���i6����Bo*���]�~1F����ޣ�^�Q����|������ӎ���G�U�w�K:�����>�/���EccQ8B��[������r���oxS^��hu�3/77�,�O��J���<d�s�XNo�T�e@U�)��]�h2�t|7
�� "��:�[q��{��b�JU�J��AW�rS�3n%�x%�-�If�В���տ��S�N]���������<H��a"3OLP �mD �Y��9�D|/#-]��"FQ}�T����8���c��^]K��T�t��B�3�Ԫa��V��2OW>O�2���f��ټ?��bܧN|^������V��Ǐ8��	�����>��۝���Y�W�����}����nX����|<xuছ�1K��������O	���t������(�"S(�����QL{�y�L���#�T��ҿ��c<�9U��y�ϱ����re��ds]�P����S�Y��6�m�C���D[�W����u��4�k��i�8i����аg�&�[.B!n�A6�������v0��P��z��^�;�̞��m�]^]� ^�&�ǁ�8���t�qkz�-y6Df#|_��n�;K1�E��&o��WI� �1��dJ��>|-�ENɐc���Q����u���}�iDV��I���礭�;Q%V���x���I����Vv�������c"��2��o��x0{�6^��[�F�7�Bar�T��U����O�AȰO��������~d�b�--����R �Ah�I��@f���z5$b���r��,���E��(�3�HqpcEj"�oxg�T�y�$���UUo���T'��ɳ�PM��j3��d[;�T-�a!S�1�0R=t�"��$j�,��
�ɦf�"Z���\K�@I,��o����[B��%�B23�q�7|��+��������v{e�Є���N��w�h�2<i�e���>�U2��� Deա���s�z-M�g̙#�+~���#�z�1��ԋ������[���B���h���?�U�!�˲)I>�3W!l�pϓ�(5�v,V[�nQk+�o�����Q���>���,"qvd|r��1+R7���W�X3G��X����;���q>5�\Jm5H�R5;�D14&���P�|Z�����&�0�&�v;l�N5(>"`9�`�I��.�NƂ>`�&?��l�7��)a������61�F�ڐ��0��0���-�ii��pr����D�u�	_�泌�3ۘ��z�����
�Dg�5g2�~Go8����&F/��"�����!������#f����OML�],z��/���$(&�CaȂ�*	n����>t�ja��M�Q�e6@-i����`L��|3����y���q�m�8�4H�)c��!j8�F�<m��7�@%7��H�-�`���5ͼm4WH*M:q���!����֕�SH\ƞ8�L�t�7_=8j$����nK�$�0s���,�~;_ޯ�Z�5L  ���;sWmN�?��1x!��>p�H��͟�V3�!$�N��t�]nCk)eh8gnm�z ����l�yҩ{E���@�wb.�8Z�fM�3'�K'���=l�Lߑ��JY��[ϐ��5���*���/�
j��Z^�X�əS���7K� Bl���IDѻ�u�n��
��K�!fg�����?���RM��I����1�e�v��X���ɻ�r=���on�g��渣i�mpX��'̫�"�b!!���RE��o��Y�9�G���U��/c��eo��H�:'���%:�'e9O�!I�����Њ���ѱ �M���'7��h������哎�!AWL�sȴA�T=!��n����!�,�Ud�{%	#��Tz)	)7�h�$�mo�5�f])ႌk*M�_Ҵ�e��e��n\�K,��|I�1C�^�5�y��
�����_�G�uW�+��<�Y[{�.on>!��s>>�ɠV�tQ��g��~�wR�B��*F�?I&�A��6]��F�JC��c��fq�����H���n����r*򫟄ﴠ }��{��}��%z�O�Bߊ���9��7�r�����"���@�#��#+U��)X������G~tB��۾��813}-�D�,����7A��N����U�'}癧�ǽsu��)a?� �������ǽ��^^�����윜�:vcҧ�'U��/���^�ٸ6�#��Zr.ߜ�H�sTBp��f�l� l���+ר��S#���k���:���2���,<_��{X&Ơ᏾�R�$�8�$5&a2Uz[�n!Ǡ�����j^��)� �C�>k�
%�ݾ��Rå�t3H�7F��k��c�íz�^�k�ۏ�Ŝ����m��&�u=ࡾ���T���'B���9��`��VB�7���+ˉU�6@�Q� ���=���7��
o3�Z������n�����X,~\p?hd�rP!1����,�\��eސ�pQn�5%�Wi��4����s�X摨v�_Ւ3iZ*�se��������Z})�~���қ�����S��k�}	b�an�P`���X���rt:�ep	{Yr��X��ͼ�&#��mw����O�f���F�აG�g1p/��,�?~��0?z�Ҍ�\Y�ci��K%c^Ҝ����F�tUNx)�����
*�dz�m��C]�d�ō�Bh�z����`]x�<��������	-�p������m��H}�3D'��X	+}i��d؇K�zɉ���὞I����`��n}��x�۹
���o�u�B�5�~��نb���tI����霻@� Dd�i2��/l�*��L��
Ƣ;aC`0�q�Wa~�j���7X))E�����W��BٿN�Ԙ����XJ�A��ÊjF��{�\�y:h�_��%I������e' S�Kp�6�&{���0���	��SZ8��/PJߕ^��\5�[ڸ@)�>�$K��o��~��(�=4�͢�wYρ�U\ErU-�1-;C�=0j?On��7���c��;���}�ҶY��BAЗy�䆄�����A�]��r���Gf���!��*�Ջ�\���(�.6������Z����[okD7rK4�����WK�AX,O�&��K� �*V��ldO(}�ER����0��½�{Щ���Y+�&z��Un�te�Z;�C����U����PeK�{5�čZЊK�+���܄���y�/Ʒ�,
�
D���C2S�02XHc���R��u��9o�E��:n�k�v_R�h��J䲃5T�3�V'�ͼ����$�ʎ�Yq�>B����A��_SF�)�rV,llӧ�������Q_1H��U4i+���nlҧ��;�#��c��c�
�J�$��^����hE�N�Guh��H����1J1(����u�3{7���WN�;��߄4�0(������vT;^��O"%V�׵�U�SG���tդr]��2W��{gV�;��g��n��*�%��A',P�r�	W|�����&3:]'u�� S��&�=��fz	��6Gon���D�U��:~�t1X8==}�l\:�w�Pl���A���b�	��V��٪�:ez���e�|`v���.�d��%+b�<l�|V�'�廬��d(�9,����v,�s�(�fm�=�Z����O�,=��i"�$��@*Q\'����PI���gMwU����239���O]	�o����U�m��kmU(��ʗ�#�l��$/�{��(�r##R��!���рo���E���K0X$GőѦ1��j��mɔ'��i8�~�����v��� <v}s�P%+�����d�Z�,l���]�Hi��������k��������Fb7�%���[�O�#�Js��*��:�l��b�4�n�eݔ�&)�h�s=/Վk�,�l�r�W<���+u�\%7oh{����L|����UJ�2���9�t��%�������\X�d��V�'ޓ���8�}��섯䋘���D����j�pO�<"��'�_b�� >y�����P��g�s����Ƌz���&�1�\j/Vl}6�|��� �*OdU�K�����^�һ9�^�����L������k���I�2��N�Xb`cJ��W�\�C��SR)��<�:w����M�61��4o��Gއ��p�(������}`7�����qM��r���o	+���U��;\ҟ��׺|\v�S�߬8߬V(�����r"���֒+�'RHx���)�U�	��=����E��l(�I�/��94��Ȑ�NPks]��rdlgg�t�|3�[tR�M�"G��Y��5+5�w��y��_|��,+��h�v3'�&{�]�8��^`��6f7���S��T�f�Iv|�"0?D�B��f��K�\_�DS��,H�U��W�=N�lڅ�>����~��YA>�O8A��z�XA��vC�#���{�*2p�p#C�Ed���������w b�XæF�����ʍ5�B���P�{(�	�K.�#�nX�;��$=�W5���iF�>h�O��	\�(_�nB��[u�c G����iT�*�����?��2����-��;w� E�;�����nŋ;www�Sܽ�w��3�L�%3���9��n6~6F��6�5�͐R��~o�'ǗZxh�,0`��������>�?tl����I�{�v'z^i��-�~*�����5}cegj��w�t��?*���1A�Ű�83�m�'w��I#�ad1a�ы5��5~w��]�߽�a�6I>�s%铃Д$���3�~����2�.Ȭ�jɤ2�;��$�I�6��DA>n>;���Ӵ��vˆ�wIq�����Z�C�>����j�N�����AT�̼��*<�0�`.���6���;>$��q��_P�9�Ȣm��ͭ�7n����\���ש��5��w�+ɚ�	DM��-�i%f�Xq4�W�_>q��%H�������N�6��0z ٯz��|�0]�CȘ~��۞?��c���� �+��)N��'����qY?���s�̲��|8�
��O���F��m���/�������n�N8��P���3�~�nFh2�v2�ʂ/����N�D�+&^��R�|ݖ	<��T�+�n&)�j��:�EM�<ƱH�<�����Z��c�k���T?׭��MX���i��̭g��-���bVLL̝���V�EyE5��G�V[�Θ����eG�mI?7�<p��m/�я?��8���� �>�L� g>�~V�?�����j,0�$Q���b��ᮊ&D�2�ڏ�ܷ|�YZ/ ]���?}���b#�{h��ˑ���N���������"�+�l��?��T"�y(��O\,f1����̈́�:���
aɗ�'�O�Y9-i�fѦ��&K���DCz���"fU�:��f��ܞ�����K;F�ьZ�L�Ҝ�բ�G����@�Yw�s�>�jJ�}+g�[�	����$��B1�|��$�5��7Ǝ|u:�]�j1f�j����y���.m2�)�>Q~�"F�%ݎ�p���OO���͕�lB'&<Tht�^4�oZ�B�_N���M_~r^^$Y(�t�tQ-4��#�<��`���^]N 5�5�}(}�I�E�ՂAt�JN��׊bZ�'v���*4��C����4}
>�xTU`���*��ւQ�PZ�k�V�S[�l�?X͈w���c�����;���10,=�N�2%_�#CYUʘ
�2(��<T���g6��c�R���M�s�0���w����ZUa��if�{�ggg�1x(��6��!I���E��Lģ&'�{Wxudk�UkU�޺��̒W��n��n|5��[6C�zTkc�\����݊m:�:�1w�%��ׄ�p�k)�J-�:��9��m�V��(�֢�'�8�?먛
"��������^��]��=��������ml�'5c-/Ӫk~wI���ԇ%��ƨ(q�'�ᱹ�=��l��O��'�H]HG���o}��V�T���M�.��p+�M}�n�A����W27*���5Uh�X�I/�Wi��=B���B����+d��2F}ʍ�O� .ҬA�f�[T|�]N��ML͋X����+����>����<�t���;�'VzOnK"�q 7�@��(�]��i�A�Π������'K���AN5I�;)�^�7�7���0'W�L����pI�6zO�	} Շ�I�VE}��T�q��w�{�e9)LwA�`u�L�P����б5�1͟H�/������32A)��d_��CW�dd/�OK��-QW���Yq�7O4K�?'�۾���wA�W��L#.����� !�^y����Q�쇸�Z���f�g>Z	�r�(åD�*m��m�Vz@H��a�&Ufj�gc�$�?�c3l7���E�mPK����pޱ10JH��Q���R�C��sΡI/4v�U�Y�@8��z�Ψ�����>v�GD7�9�S�b�V�3����EDt�e�+$��BA6����WJfPw�ŝ�q�79pT� �d�^��V���̖76����Γ��D��H� <axs���""��.h4�M�`� T����ϻV<���4y�YN���t�׋bOJq ��+�p�~M�*V����+�^ӺG#|�uP�ZVVó�70�G��㐦LPvXe!=$��xq/�z)a]=����m��EI?x	��RC�F��C�E؜m������ؼG)x'�v[���$������ɵ���TʘiJ��X��+��d/�l6�t�Ro���ΜWD�T� ��T_;,Bn���v���G��fȍiƮ	����q��b�o(�ڌD�'�v�1�&�8]~UY'sr*�V�ԺU,�wsO�����s+��G����F���֡K#+g= ��8g���X.�/͔0X���v�~%)J���b	�YH�S�D��B�	��L~�V�<�b��0ɟ����]�.L~�A����*R��#�Bq�Ԁ�к�3&�b�P�Ee�0r_�y���������o�"U�j��'#�YF�K:S��:E5�1$��e5����4���͌Q��,��9�����5�&�9��ť���w�	ܖ��D�S|`�[�i�^`���{��ʋ�ZY�բ�"�s~��s�A5��By�ߗ����[2lȠ�MI�K>��9���<���X�D��U|�����J�ƿf����&��*Z.��?W�4�T�!�PEz��n|���ŐG|Vy�@�&}M\	����W�K]	ھ��Y��!��0Ox)����S�d�r��/�KKO�4ag��8FAH�\�I��>=hsu�PK�������|��e�S@��Z����;[%�}�U	ބ<	Jn��0��B	����f�n&�;�vd&FT1oE�e������_i�*���l�-�����l�=�[��ַ���Da3�mfw[�hu��"e@�V�ş������P$��M����ҽ�M)t��ɳ��Q��S���) �h�j?s���ױa�Cx�+�bb�Pv�!2�o��b�4�;SH��(��\ ������W+������8���885�������)/�v�x�����PpcH�1*q�M�Q�*C��JV���1�A�2j ����碉�o�仼5hd+��k豟sc-e�[����~~A�<�Ċ��:]��8��e�%:s�4����+������6d�e�f>E��u��[qk);�pm��x�6
x>-g�4{z�4"�s	���|��(��
a|�f��H0�W�����{�,�� �x;:�ggg)W�����LOO�	��e�r�ГJ~>~I����,�锚�Q(2@��s�"�V�6��z�%[<��9��>N��P�RZrRX���
�L�7���2Lǻ�d�|�*\�?nOY�a�I}ϑ	*K�k��V��ϔ�+�a@(�pY �`�M�d�CN������Y��XY?�s!�߲�2N	SX<��"e\hJ�������b�֨�}�����sX(%c*i�����L�M�i4 IСHOɫ/LL�>@.c��D��!ڸow��e̬&��L����-�ǅ�H��}�e�m�͌#8�?��d���H G��
���	z+$߳�zy�#6K�=���3�v��$vvv��sGYk�����ٞO�4o(Ұi�g;����p�:�l-U�Jb�^����"�(�siBq�%�<
^�n��r�l�N�Z�$�e��t����j���<ȅ�-����.���,�!:\���9����(�o�p���*����ꗚ3����\�$s�/Nu]��d��\/!n��o�/	KW�i@2e��)�x��EmG�x�h8�X/Rh����I̤D��u ~+�O�H��0��t�/��W�4aQk�O����H�5��]��β̠x��3�!�����@�U��^
���Z&��f��I����0_#P���������	tOM繲�~VF�/��H���Ł��V1�T㇅�D�e�>�V��-JԚ���z���T�k֮�8]��͑}e0XS��F�����س��\6�~�Mx�Z%ڤU�N����6ď��T�ē���Rݼ~�q2�C#�:SDh$���l��A���[��ݩ����`�r��3rӠfD:Rq��.8`!�g�r�r5�=&�U�[$c,x��},���L���\�AA$�^�Y�뗑�\�kĊ�?��O��?�vGHfu���<�z�Y�w�>�������D!{w"��3��]�#U��`� c5~�ȁ-d1���܄4�������k���4�{��5�{xn�Fi}KW�G�.�LB�|����O�����>e�	{��MQ�Φ�ҩ����ܘ���'�Ёr����������}K�䜢Ф�_���ЎL�4�hw�`T��S����8FZ4>&^�ɹ�*Q����{8����v��*�*y5
9PX��I�,���L.�]��A�'A�\��B�g|c�0^%s�����S;��F��K���e�"�\�+�D>�Y�&�1؎��ʇ�Wڗ�?��ie��>�M%y���	�������Oeu���h�6��-�X����&ֽ3��|�>��# -��ypԈ��d�������8^��/��駬� bTC5d,���V*؉��{vYr�!T���P��J��x��=�0��Q��h-����R���`ٕ��p��e��'��m�W�=龍|n!a�����wf�N��FyQ�����B�H����#����X�v;��4rL�s���N"�q#4=S ��zj�"WO���ki���3�M?����ܝ��aM��>
'��D�ј���a������X��?�ʒO��Z2��<�D��FiմRs��O��Ef���,�OQ����>�BSE��ס:r�pd*.&p�̲%X0��΅�Ӊ�T��6>��gH�J��y�'����Yb��R�%|������!�;Ӯ�юfûg��%J�H|[�G-"Aِ�0>T0%����Ȱ����8����CAD���w8Oն��=&F�U-�����τ	�?�K��UW�i�>Bg_ۨo�k�a�
qy�;�	b˷���ST��"�fĕ��r-��vN;c�_r�{yB�.�.h����q���d�k+#��R"~9Jǰ;Z58�
���Y����f��ڀ>��&�M������|����,�c���a�9�nWE2��K���$�K�����e)�;���TF���,E��7�v�h	����{q�E���nإv٥�9HUC�vQav~�o��o���5K7�*^����!�W=�����4��#�Z�'���|�(�e�3�,X�5�&��9��p�X�G�;o`��6'�^�O�6if,��4ØOe��i��!|P��s�V?+��
7���B[�v�W��i���<�T�@����>��:!PF��=��i�k�2w��R^����V!���O�VY�s�������.�PL�gEs�h�tw^��ٶg@|ˌN�(��K����dϋ��ǁ���%�W�t������:�._��(Fqs}?w�[g�^H&f�O�[����5��%���%
���ar
�Ŭ ���g�V�3���R��"ٱqp4S �7X"�f鷯��w[��U��|8?A�[������.G]h9��E��7���c��{��^� �X�0 'Q��$���rk��[X$ٿ.�qvx(!�V�~g A]mm�����F����}�m�(C��Ԅ�ѣR�N�X�Nk�C��uB����P��p*���X�@��R��g��"[�-�����>f�B�g3i�-lUKxal�.歝�T����@�7��z��;_�I��Gq�X��S�e,��۷h�^'���,,��#ۦ,VE�_���x�ͮ�F�Bi�������
�'	� %{6�g3�%f'�;�����k�XkC�1T��O T����{==$�%a��F�_�z��]�j��LԦ3Y�	�I�%ʖM�|����޿��W�8���Ic��-K���V��Ϲ����7d4�Q?��fg����z��B�I1p>@���l��r����̖h�����˶��2��3!������w���_�η7�H��kM%�6t	��@"�W��M��Ժ�ʖ����K�n�����
���t�,	�\-}�?��sICW��}��(3�sYo��:����&
�Y5Z)�a1q5��*g�J�,)ٮ㻳dHZYx:��U��xC<Os\�Nv�/[m;P=7|=�����e���w�/�~~9�~3`5psK�����Tf��v"�쩾��!O"��2k��]��(о`��N@�b���������y�#�^���NJc�ؘX��cƒ��R��Kn�9�HhP{{{S���^A���u4��6�W����E��5,]�m��|㾤��dV?+�-��.��/Hz4AJj8�Aᡮ�I�ӯj�P������`]~'��͊d˫����s���֯�,oŖ������I*w���jc(�YߝÜ���j�}jʭ������:`��n^��oR-#�ҁ)h��j=W蹴ç�C��κ�ԇS������<��X;<,:_�c��M��څ����\VT�U�ަ*Td���fU����Rs���.��^z#�2���I7�,�Fs���0�ѩ�u&x��e���@�7=��K�\���PD\M�QYW�މ	9A��/��q=�����|����@�a�06>>�O��	��L	6��5�ft<i4�%+�t�WZJar�D����/�.�Ӏ]��a�x,��R�KR1������dvD9��{�{�b7PK|ފS���<*�&��?%}�+�nys%�2�,�(�a,z .��[���.���-q�T��8�����쁍(�U��#�Dt4���/��-V�6�-�Sf� �R�ת�(�h��yY	I�C̯d͖l[�wߐ�}U@+X ��h	FDF��{7�ws���+���鬝���[o�����?Bg����CG�|kɽgXU�٧o�V��˒���j�����2q�c�.��ոȞ�ē6�~L82 �=������,,�{�C��mr��F)Q�=8i:���@�i�`��N�[��^qBdPN�9�b��Қ��_��.o����<�
s`��t���ʕ�FZ��QY��!��y\m�;Q�!:Ȥ�Z:v����<Wb����~��笋�=n�)2�)����xl<_E��K]tj��YA�H(�V���G)�,�LQA`ˇ��R��í.Ǿ.��*$�]O��0\��*6��ۨ���*{��yif��_�F��Z?�=����B�����)�Ｒ�F��"�h�{D� >�C&�r�]�����%,'�P��f��� VnS+:Ş=ňˬ�}t5�YP������������e�<^���#�h�����+��d�?��M2EF�I��s��C~|�zD�e�"���L���wN��&@f�m`MnLf.7�W,�o���Վ���������F��~b��)%t�*l��'��U�0����0�Vt[���ew1����%J���M�0:]�}g����7Eab��hƙ�J4sN�QL:S��ʔ���}�����;���F����r�'�~g,:�5����"�V�1I�q��)�kң��Hǈ�@,����T�9���I��e2������rǽJf�X{Y� �h|'Y<`z&	EB���.ϿE#<��y{G`��M;�e�����}u$=����^�ނ�����Hk�/Ɖ��Y��f\(-�)�HB��hvw_��عU���<�ؤV ttps�n����z��s�8���ƭ�D�l���nuuӫ��'+U�C��V�D�ПN$UjQ�77��|[Q��l���2�y/3�8{�zz�¢^�g�j��a>����4��F4- ��W�6iU]�E�Zw�6���i�A�<��KI�ڰ7`.�PE�Y*jiI4����� R�A����sv8��w��$����pc���NoY����%�)�w@��Cȳ*��S��;��4�9*٦�w���a�� �296���l�����/���g�E4<(C����}^�V>����M?H$��/���]�gx��zV�z{�np��[N,��-ZNMV����L/���2{��X�����o����z�ۚZ��/9���W琧�X����sE3Je��$Hr��:2j��Va� Vt���z�'-6�R�F}� `S~� W�5�0������c�g��s���r�~tq�F���8��X�e�>���b5���]�PNY�I����F��NO����|�����#����X��`G�����p|z��g�P��O��K��,�,��+�~8�����+��ΝoW��.�x��JԮ����$rp$R�ZU��:QCO���&3�8O�b���*��m2��<qpy]��,��!�l˙�LCC����t	�%�����Vy�ݟ弌LL���?��G��	��wh<��G�qYu�!1�"K�7 �7����9(η�,*Q ܰR8c�f�l�
��_����8A�v�,Vtl�Ř��d�a��Y�o)Ɖ#Io������ 
�zd�oT@Ѯ�@֛T��ʜ!R�>V[�q28c���}�T��@��'�?�j�ff�H��K�^��'Uj�4�UUeLȎc8���t��~�3�h��'����B���0���g'i�R�oJiӌ͔T�T�	�X��(ƕ����Y��6-G��*2���-�h;2�#����.��&!�2�^\���=��{�����j�	3�HSn���<7�%�:�uZ��ύ�P��B{oDC�Y[Z�:8�vZ'\yU�9	&��de�� ������ʜ�Vd�`F�ci,#M�(-e×�#l3Ŕ~l�I�&���G�}G�gJ3�˭�Xg��]=d�v�ғ�e�T��tT�!�ML+3�B�"�`F��v�Uwqi�fz;Fo�*3;[\fԄ���-vEq����-ަE4w�_;��L�� �sbr�HVx�io%q&d��By���a 7��|`4�A�VO� =;�<U]7ܯG�]�SjkcC���T�b6�b���E �v�-�;ᚺ����,����($��-��,=��
����-k��,]�CQ��Mkm~5⢴��*�����p�i�A�s%�q �����$����;R�i��E�Y�VS$x60)n���d�`�;��{s}��{?=*��b
]>|$�8m���l/��-}��x��W��wl�/..��Y���D��#�U=�gi��Y�`��,��}��o�xa������`#G����:\��gd)�*���.��*.I5PG���7s�GV��G����� }!�)uL�����;�U����H����X}���Ł��=^����Bne����������9�u�uLB:6�ē��
�B�[���&|6���Z�6׈��R�P]��w�֩�]�%9O��~���4�g�j��®%����BSs( �~�*+x�Wed��s�֕�!�5�	@+W�t#D��?�͇n�=�{]!�����ߥ�B��B7�/B�Q�B6���'Ζ��x�d��H͖�ײ� �8U<Z*k�p�z�_ �.�Įl�|R���7X��m.w�4��8L�m�����nt��ݑ�ib�AIA�%
{qa�jjjx(�|nѩ�O0)�u���1�@�ؽÛ�
ܧ�D�@��P�?��|0m~P�y��;>;���H�4�����>DQ��޶>�I޷�^�1����]�r�������_��ƀOT�n�f� �*P�"��Xm��a��PQ|FڐrnW�����͋ڏW��#��읺Op�������_+���{�k;E�)�N�s�<��f��"�<&�sd�,Hk�<vO/T��$�(�򠜞�����y��2H�ea40�]7��	�r�)"�����"C����?̐�oI"��H��X����N�kQ����,o||\�B�\s��O{�Mv���u���4<�����GՂI��������K��Q8��[z ����B� ��7��׷-����s[�ic33j�20�8�w�w��Xq{��L��<c`pޒ�3�1�0@>��{��=W�����0ͦ/���߶.������o��E���z���<S�,�h9�8n�n�n2��c�O�+q�[��R�Z�B�S�9�BQ�v���T��e�.Ԝ�?O��z�#��F�^7�u`k���Z���U7����j�����,�!=;{�N��gz�nGeކ]}#`��:5b�Hljkc������5��|j���z��cy��(<ׯͽ*�������_��`����z�G����.�F����șs'��'Z�n�KͰcE�'H�W7tv��>��x]�0#��*~L(*P'�O}����v�%��Cb�����1v���`���j�+#��Q�~��&<�t��*�G�V�� S������Bܦt���Y�܃P��,Y�My��@��ŭL��@`���9��fۃ���^X?1� M���	�b�aqc92�߿��O�o`��QcCO��0���>�����-����R��h���������'&��>����\*��B������ǲ�o�o�F�����H�1=��MG���Y����A^]�{t�c���7���S�䊝������/��ۜ���Z�W�y��w��E�N���x�e�ic!EG�!����vz���/�Hk�AW�m�=E"\�P�����q�D��]�������?=�_/�\��a#|8V{]�ߧ�/����)�z�%��F��v��E�g���9sq'�縹�o���_�������9uey���9�2���qin:W���0�I���ˈ�ʩ! ZX�g�_����pY�� `bݪ���n�����}k�S4�8��5�6�C�X�ؼ�t�� ȐT��:���{�9#��T�9����Y�(5�)�]T�$��	����a������9XǨf��/o��'�����p�����)��"�����ҳ��xM�K8;?G"��!����Ifq�9��B"(�4�����WbD(z��P�`����%L��m�l��P�Y�S����f���`��[!o����$�{.@髻���`=;��� �VEk��vF�Ix�u�(����\[䌅X�M$y�N�u��S����z��嗶3/<��eHbX�\��U}�;]����Vw���Q9�454L|}���S)c�&��[���m2����;�ӛ��j�ܭ.�|:=�17�Ij)+]�X��y2������:f�-�F�.�5Tl�$�/� d#�aT��a���n��>��Q<z��"��S����KTD1����x;p��q�X���`�}�Ǯd��1F��/����3
!#I �/s�X?:��K��l�"����]�|��n_����+ǭ�B���d*"�]u:
�ֶ{q����4�����,�9�u�XŇ�II'��D�K����	����=�u^M;�g�\ߒ�r����=N�N;�7�;��V�^ɲ��J{J����`��'�||GǙ�j���J]�l|V�bKQb�r����`A/oI/��u��9Wh\�}�cĠ4)�j��C8W�Fo,-l����^}����u������y6�\�ް;�_p'2W��o���R��3��F�2���S�Ý.���l`j�u��O�����a��N�9�����?�P�P�6�0l�1���1X��>�?0k��2Ŗ-��,e���0U�U�hi�n=]�ۤ8�ʚIcK�֖�A�p/w�J�A��y�m��c�>���@�$׾Lābɿ��;�*�*���HH���_�/�jz�s���{�6/p�}�5����GkÍ3���t�N��F{��>Htۜ��@q/�������[�^?���<]��vݠ�c67cYO�F�T�z�-�0�L��%��:CP?�r����,��U5�������sm�s�"���B�����@>c��v0l<�H�,�nU%�Q�m�CXN;Tf"/���a��U�2�(�KFU�]C�bL��v%0L�i�|�+�
m6<^�]��4=g��u�j�D�����7���*hOM�\���-IlͲn`g8���r��p�@(�8��s����<�*[>��/,�S��䘅�{�����=�E�=-	x�}�������(�,�U	�by�g�%�b憡��Щ��
$]�1Ԡ�����rI^�@BO���#,�o�qY_ �:��]1�%���}��V]���/��1h�D�h ���92\�g\#����ttb�"Uす�gUL2S�>�`���44*�>�k>hˀ@�_*�3˙?�����Y�U���׶��..P0�("���:�^�eY� �d/J8��G�Yn�W"OOO7����?�m~�#y&���e`-Yl��"�e�J�@0%ˆ륖
^}�y�W��L������������3���������\���ja��-�V����p#I�T�t��'���G���~�W������8��e��K�O!��}2Q$��y
ټC�f��Qv-QhAmm_WϹ ~����l���xB���PY�U�����!_-K�M���O��b_��P���.b���C�\�zJ��{<Q�4,��×*�j�rwr��lk5I���l�&���hn^�T!� E�%kh �?`;�9���1H��*'(L,-#&�u�.%��)婒eB����^�5;�b=������:f��++�h6u���bq��u��q�x]�����s�wGw^����{�lC����T��Gqa:>o�~I [���[���p�6���%4�+$���=va���:s���!���"!h��m,�@�8�'?���N��z\��b�m�#O�O��;#�D�� �%� ^a�`"X�z�Ћx삳����7O�����:�B���_c;ÔQ���k��٬b{w�%����NCj����g�Xi��>����a�;�̡!qh���^���'w� �C>s��h�Y���`Y�ܳ��eE����))�x�ϐ��t��Ƭ�]��a�.�B��ߍoX��;I#����������&Iҡ��қ�.�։��j�*���S�g�Vo�Aw��Cx�Dx��Q�=�ŒZ��9�z�O���}�f����ܩ�tu*�x(ԎY	2�����!�"�pa,1�39:��
�v��͍��D!�B�������$��Ѝ����ښ�
�Eb��d������$Yф%1����@	��:]a�u���5��Yiv���3�6E$/�b��/3#�kK(o'+�)[�Y�#s�1qu�/r�D���]���dFw�s�m��Eۮ�(�(
�gͥ[����c�u����nF�bҐ��F̥�Ʒe�o2��"Z"�e�.�58�֛�LN ���њ9{�o�"?Sҥ�9ت*����åk��$���s㡤k�n��5�h�~`�4�E�'��΂�N\�C�7}��e۰2�j;/d�Mu��[��ѩ����C��a��l&<�o�nq8�Q��R��rm�x:{4T�8�.�w�u·,>#������O�sg��|�|��6{S�z���W!�̨��QH[�N��ZЮY��9%�/�}c��N��\��eL	q��ڤ��sL��/F%7&�9�#U����s�0�Kp���<��~��c}�7߻J{z�ș�0&��>�пg���P�M%o	\��_�a)�Q^Z�[�xt��`��9�+���y�j冟~FW��T��������Č^g�Yx �`OV�BVT����|� �Qc1�j�2E.G�ڽ�D�ݑ�eW+C=�u`�7OlYJ���m�\"y� �\�qOOZ�Zy4���X�V���q.��������&'J��bݥ�˝�r�$�H��a���W�h�q����}�5Ѫ;5��D`v�-�(�9S�,ҋD����8md���94a:cL5k�v#hr���	�lY�(z����$�X��zJ�}kl�mY۱FgQrRxC'�i�j�}�k�7�#1}X�-k[���$����S?����8m�c�P쳖�/�rE�hE�z0�`Qΐe�T �jq��bbu����S�pn1�y��es����ï���,��6��l�4�u�±޹<���k�	�<�"��(�8������7s ������(���,�B:�Z�V��8��ā;��/
g]�\�	�=�Z�nT���9ު��3��2E��XQ����
S]���ܨ�sP=���`�2�����Fw�!�h�6�Ro�su��4 +��cw�V��WWG��:Gc�ː�t ���˛��	���?2�n��k�ٶy$�g.����^B�F�T,�I ���6�����+Q ��G��(���odn%�Ⱥw;&�c�S�����˥�!�wq߲�t@V2���-�9�h�3���3��`nY�g�wy����m��$]��wN��X�b�_���/�-1p5�#3�8��mw�PӒ?%ٿڍ�!V$�,)��iAͩ�FW���X��	��g���r�(�"1�tvO�4�N�sH��Z�2&�bY�Ml�\p��8�A�w�>�o� *�I�"�8�_M�#������&<�����>S&�4��'������ݹ\^dbno%�!h����� 7�#]�W�L��a��P�pH��0��\�d�m[_'���Z����i�ZH�[91""�O��B' ��gA��O�=���Z�/�L�t�q�xH�������E+��j[%:��gn=�(�Z�T�Um*��:z�p��8�cpH�m�ĀY���/ұq!|]�n�T�u:c�~�(�4��1I��{�o�b"f^=�lEbH�U�7�����"�nk� �tj,P�W�x�+�������D�(U�
i���9x�q_&=&�U���j��+�p��ɅM�i��!��LW�Ѡ�N��])���f�e�@�7�І!Idp_�L'
���1�W^o��Yy��e�m���?��>j����ESR�$����Exu�,�pf���^X321]-�t'0�|��!�q̝W��9o#X���g��w�NNƖ�S�s�s����_��E��4�+�� � F��8YU�ZSS�b��Udʟ�!p'�	��B���jtk�liפ�3Y�a)��Q�ȑ���)���l�P�e#�s|1ݥv�|(���pd˭��C�ף4e)c�����jz�������ݽ��{	���2[?	����)rw��ާ ��q�%�.�ŞcCگ��R�z5�Uj��#S�u��΁Uj�MZ�#R�������\�ǡ)OO�!@G�eu^6����P>.�"��
-����R^��_��* ��h�v&��N�3�r���ڍ����{�C��^�<�k���p���2ؕ��~D4I{J�� )��aL�V�}'G���#���O�05��6����c���Q�ϙx{g�U��ࠚ[Z�� D�K�I\-Z�_�Ga���
)��"8��.\w�{"5���!R��_�6����ҭw=�N:�'=8�F���}�����\����'������	������s��D�P�SR*XQ"K�;����.�+�y�T������E�UO}����[�����[�[�O�?�
�M���d�R� T	y�+�8�j6�-�^��j�CT�H(7�������Po\��f>��[of�GBL��Mră7�.��sR�u=Wi���	�K'�Q���C�%��Yh�����,��w('���~���r���EɧO����(32�V�
]o�J6��{� ��Um�����?f���]���nұ!vTSB���P�^���s\�����}�p�"�>ܾ���m����@�g��>��P_����=V�'w�M���7���lK�X�ؙ��J?�f5��.�m�2n`�͐r���89���DK�պN�ء����~{�BOe���k���u�9d��cn��%�㖍g[�9��49�ȿKK񃻻�QQQ廤�=5~�C}��Y!Rr�h���3V�[��͎k���${^݀�Rp����([52Q�j���?T-X[��w�,�"��=���dEZ\\���0��K�i1�����I���>�Wۢ����0U�D�j3!�3�>e�l<�B%W�v�~	�D\>��ַ��Z�JϪk�@Ғ[G�i{��⒝���ԖG�Z����W��(7QK‾q�
�ȡW�.=k����QN��ƞ�Ƿ2��g&1�w�ѯX� ��:O�w
���	qފ
x�l�
Ƞz���^d�;�U��r��R�{���Ln���};����tz�j��wf3=w9}� [:;'655eEc��gffBD"�@���8�(�Ѹ\64�UЋ��ަn��u��_8_4觋�=�;�C� $HL+&P�{�KJ������6�,t���}%�#a#��\��i��@�G�����U�5��V�;���'�/��1�F��O���0~�u�]�-@�!C��M�A��=7�AUĎ���&$���H�DH��%��EJu�'E���hm��� b��n��\g�r!��2B�6��b�J%�H�X%�X�Y/iUlE1I����(�qm�A�O�\�3�b4��nUpݔ�GzؖK����� b�2 z�i����^�i�$QJ�.A�R�*��Lc���qf�[�F�j�Q�TH�A�n�U�c�C����	���)�0��P`:u���t�v	i����b�R�E�Ӓf����}X�����4�X�*JlW�.�0-��d�_d}}����#�x�	}�Qj��-g��%��o�[���C����2t��^-ځ�ǃ�-��D��4M\�ʄ	�]�ڨPkT�T���Iӈ��1�� {_��:��"M�:��R������v��=3�b4��	���rU�@��#��h��y��@;Ƕm�l��q1	T*ayyY�.ʀ��OS\ۄ�v���'
#�E�eI�0���׫���T*Ah��s�q0��!���:����B}�h�PVȃ�����l�a`����^����ԛ�\�pnFQ?����o��?����q��M;sĉ$#l�D�*ި�.j5����dr���o|���2á��Yaw�F�R�Zj`U��kgwHeH�^%
�*��j���ʏR^� ����T*�!X*[�u���������n �R)���O���[���`yyY	(���.+++DQDw�W�7)%�dk�:�e�x'1�SƮ9XV��q��0���E�\�U�LS����U$�{��#�u��Ϲ諸U�o��G�D�E�E���3�ʱ�1��$���$�^ل&�&�"@6Y8�d0�ăh�I&�c�2,�{L�"m��~UU��>O�ۗ4�T]�
� |4ϭ��s����}F֓�#Z->�+��e�֤���zY��EI��k�Z�^��0�p]�;w�G?�	��/}�K�~�"wn�&�)�i�c�ʏ�7=B�R�0(�H�L#k�?B&�c	���7�Z	��m֏��?�c,L��0A�HbI��yP�F��D�S��K鯞8A�QG�U�ya�4}�q.��aN�(��u�I�w�!�t����ȉ�8�J�G���p���40=H5A���[�6#)�	�j�1�ZI���z]ͤ2��޻Gݟ��H�n"�4U�2ɖnt/F)RJD����f*���x<ƭV�Tk���U.5�ط�!��O��.}�W?����q��]�F*��G`�T*�Iİ��^�id��\?WG!�n��O�������'>�������m���$XB>�U��	`96q�0�#66_�0>��#����kTj5Z��X�	P��.&�_������&.\��T�	'gΜ����� �kд1�uj����]\���5^z�%�߿��%�vU���l6����������ɣ�>*���0�a�!V���;C)C��+�A
��x����/�������	���p���u��Y�k �m�L%�h�1��0O���((�I�`}�{�GKV��y�3�4��#N�<�L-�j5���}~%���eBO�-􆋬�B@G����r��I����nﳶ����"��V^w�m[	Ogan11W���J�QC��2T����&v�S]~�g/�η��J�?%'��B2hu	{�c��wh��sok���e�c�� ���6�qH���N�����9���Z��NP�I3
���F˶��gϞe4�7�8?u�~]MRk�����P��y��wI��Sm#!��1
�DA��)�s'wn�18�2F׭�oY,/���ɂ����AL
� L�D���2Q�k?f��o1d��8��WU����*�7_ckg�ᨏ_�9~�87o��kIE�0}b��a��eZD���BR$/��"պ�aܼy��/�b�)�x�iC旚[��؂PJ���?��?�Fw�E}q1��JS���}��a� �a<�a�ק<<%�[���1���M���>�0J�Z��ܺu��}���0vk	�2��lp��\�r�o����B��;ɘ4M�Pi�����2���S�c�;V�IV�W�� R*��f�cǎ����o����eww����4�ƃ���vH#�(ngo�V�E��֔��:=V��4M� ȣ;=���\�É9!�c#b���_�9�u�V��a����2��I�6�iX�Q̉��p �6���t��F��82�	v���ؘ�E�WM�K�����gz��Q���̻ex!)�L0=��8h��dt�8Qw%��!z5�{w�x�w�8w��u�kN�P����y�p�{׮���!��2�0D&	�e���`��J1
9���� �˰iz>{w��̨�	�шz}� �#N?����.B*
�h4�G���cG�qC�a��!v�F�v��k��`���O���2Mj5���}<����$�%/.����-�����V�E�9�p<���3�;-^|���9�����C��0BP�}���XXX��HI!�j[T���R�$������Ǹw��/���w9~�,����I���p��9��ܾs��AhJ�~ �6��v�� ���H1<�B	��TeA
HD69]�}�fD� �b,�����W���A�94��*X��Ƶd�V�0��Fܹs��8�>��I��4�sz�Ƈ�oߧV���UfZ�R�!�l���Kc��G7>���$���l�ߺO(G���,L��a�)�r�������GW����]���uKU�ۭ��q�zD��iS��Y=��ضK�a2��K������������v�o��t9��
g_}����g+�z=�D��秋��&RT=�,�$�0T�F�������4���9d0���+�� &��D��	�_���[,--������I��n��1 ��K��,��F�US�!�>�i����:[�c���K���a���UH�'��,�y�j��e�� ���_�3�}H��� �0�"bէ+@�b`H�Ȕ�D!�4b�s���2?��x&���&�%	��1̔4U����/h�]n߹A��2�p�����$2&��B�����1�G�������.�N�I��ģ�������txU�URo���wh��BQ=�]����4���w�JBFq����I�ʢ�:�,�J�cm�8?��2Y�ۘ{�昛���'q�):`�)],�Cn��(���XY�N��ad�Wf���Tƪ�t��F�.����m3GHT�EA0���f����z������j��=��m`��,4�$��4I��$���H�È$N1��t8y�,���"���[�ܡ}0��X^�(6�1�tq�
�b���G]�$ �F��T��>�h4bgo)^9�*����%��N�K%$�Ķ�<l�!�$!����7	�1�q�51��Li�����dnn�n����6RʼH�����y9(�1a4D	�a�Ѩ�0b���[��s�c�YB�D�iILK�7n��f���-��:��~���$ID�D�1$���k�쑪�I�5���|R��xj�
X��EE=T���j�
�_�%<� RSҬU�l�A�mJ\��6!�c��׳�*��K��v��yY.����Q`�:s|�w�k�^f��݃��P`ul�Ǳ�Xf��iT�z��5�2����D%�eR�UU�!�ٕ�벾���ٗY\^�Дǜ�!����\u��J�e4��u{�j5�{�.��ַ�F�͸B ����8�1�(P�L�ƶܼ`x��/�T]N��b�)q2fo�>�/�´���R�T��eY�|�q�`����p�K?���:T�l��2��EF7�lLS��	Q��:MS�ՠ(#Q�K�$���01-A'��,�[3����<**��:�T󾑒�RI�][t����矪� �ǲ��Yẖ�����0"�b�PҘ[B
��p��۩0����`��L�ڜ���a����q�iݧ�8�A8HeB��!�z}u�۶M��Y�'���n�ĊG3X]=�������ͫխV������9??�A��@ɣ�贈a�:��`6F�7�礔�Z-�x�HF��׿2��pH�����ܼy�S��8P|�̉ͯ�ܕ�ٵ�<�����5��2U�XH�8�ÀJ�J���v,�z��(�NZv�T-<�i
Q4"�TVP�{�4lR�湕�|i��B���Klݾ����9�c�峸F��[}l���m�!�2?�Z������>O�V'�$����%G���s�4�sj�H1����{�߻����4j>�c2�P��g��kS��H���TB�|N���1++6+++�޿��8��ѣGsy�;w��.+++�;w�q�
U�6ۖK�L,K2���-s�����t:��y� �s�������n��ƧO]��u�~oĹ��z�a�H��:nN��l[}�˗/�^W�{}nݺ����HŘ�*V��ނ8���k9yZ��:�f�X3��X���F���͛ԫ1/\��n������S~����&�pY\XQ�f���쯔�P���z$���>���5VWW9v�����4}��6�v;�^����
���[ �Y�e�Z�R�Jƣ�h(f���D��&Q����N���S�n�z��F�dIν�]�����v�
A(���x������aܦ��c�����>��D��~�j�Ā�Ԛ��~������f4R�`0ȧ�i#y؀�X��:�Mm�L,JPmԱ��u�$I�����3�>��~�ߔ�����,/]�$/_�,/^�(�(�:��>�}�������[��ߺ,��w�ȗ_{]�˷ORNl�k׾��s��/|��W����߻��z����oO�3=.� �j������<	^{�?j4���������;�v��Y}��B�[�7����"��Z��'������t9�14EG��U�xAzk6ڤ��3��Y�O��6��!�Φ��bW����IF=.tw@�Z��ޫg�O7n�CWpA�0��hFГB���*	�XtΦ�N�1��Cu��8.�`4�L�rt����?K���9-�i�)� ��/Ӈ�\�"?��ʳ��u�u�i��<�@��|�~|Ys�'��5����܇�vv��L�T�6I<y�X�h4Ĕ)�2cF!�����c��2�L�p�ö��5Mϓ<���3�?I7ߓB��گ�$݅O}�i��+iB�WB���F�C����_��ѓF�����ӂ�y�'���:oQ���Mjp��U���d�b��`�w���+���(s=����"s�(vk�y�>.f�`,��F����5-B��M�T4�	C���tiL�=t]G'�tޢ,xރ�f��`�t�g13-�i��Ρξ�Y�z��2PJfY3�����,0����nPj��0m&�noH�H�p�d%�dE	�Wͅ��3m0:��=�A���:�C��&Cj�Z.SV�:�h]�g��vzu�5�_Z�h-��0J���Plڟ��	�qNd�|�2�� ���J�d0��<&��.���3m0Z�R��U=ֈ�z���U�?�ӧOO|�(��̴��n<}E��Sh�kOw ���o��Ǆ�uc�4�03���nY6f��W���M]�Ų,�޽K0����z�k��;-����Lk�l�n���{/��8I��\qt�N�q��Fy߰���}�����!�b�0±l<�x�^�4A0������Z�D��uϗO�.�tv���t���u<K��	S��)e����_�%e�Q�r�3m0�J�P��8U�$�om4zz�$�O��h��`&�z�^�����VY�i���1ד�'M��G�>z��iF��$�j]u]���ݯ�փ\�xTO�i��a��O<7�	A-+�/h�j�}�a�M�,�+�̴�茫�*�C�ȅ�ҒjZ�p1�>���6�l���~��َI�q\�$I҈2*I��*91%O6-��'yB���Q�y�s��he\��|ӆ�7��Tٲ�z���T�CZ,uLf�`tۇ*z�vQ��LL�3�Sa\��|x�DYT�� �i�LGI �j� �0�J/h�E'��q����J~��	�Cв����E�0�8cjҘ��G��?a��>�a����wp���ӥ��Q�!�3}�h����=�Q�$���B�R��Wq]�4��a�ӂ�6-������u�Hk=��6~Mݘ�|�L(�W;�e7�۶��6�b�g�x8���`&�^����j��Xf�,�7��O��&��Sa�(�L[�z�f<s���|tr��I�tY�ƓEc�Ʋ�\��i�B�ϭ�8e��E����3m0��q�����=_d��碈��է���h�vL�x�������L'���T�yQ�l8����H5����N|}���OZ�L��>j��m�Ξ�SD,˿(J�=�a&�ZM���ɢ�#�25t�u�i����I� �^����2�h��8��L�4(t>7�	a8�Uc����� yBM����Q<jd��L��ԽBOÇ�b�_���)NK�&c�78=u{i��#���&���OSY f�`t-GJ���j���H����2	�3m0�b�ia�-֏�c%�����ۍ�m�p��ɈJ�"�4������������Y����+˼x�%���Q�k�A�Z����f���n{�k���s��ܱ�<�k�{��<	f������5N��N�&��8^�z���_=}�4������������f)kmllP��B��/|�Ry̜�H)���R޾}[�axOX&�mq��}�%ʕ���u��666�p��i��o"��:�u�A.�����7���JS�x\�ԕ4�|�0�Vw���2��VJY.BGb[[[�qL��accୌ#3����H����}��$�ˉafN)�Y���E��u����V��S��8{��gΐ�db�]JyU�2Ǖ+W���G���\�t��p���oI)e�2�cY�'~)��R&��������ŋ'�q>5��W�نJ��y    IEND�B`�PK   �x�VLp       jsons/user_defined.json�X�o�F�W�?۫����v��zIZH+������UbS�4�"����9z��HH����켙��%ꞗ>��V�o��}QV>���oߴe]�J(��]e��mt���뗛��_�X���OF��G�u�Zx\���?��3.�~E���_��8*s\�$d��,qF�D8���@�����k����u�U׬��X&�uM�춁�b��t��dY=�eYM����^�j�8)��"}�L6F�e��dwmV?��4\k�E��̪*�Za�4�wM���u[��^���3b$�&�	Pf�S�*��np�k��4����<ZǇ�� :'��b�%�TY��H��o�ӣ� %Z�1S�H�8� ��:���#��0�ɜJ`:�=J ��ql���6ŗ�$��>�L���FHwێ|*T�j�o�r�{}�(�>�o{v:ͼ�%6�������(���,1\�D�g�|�-��e�CZ���R�Z�5��<�g%�Q�A��jA,���ߴ��K�����#Ty�mw*��<Y��q_�����l,��5���y���)�"�,T�򂦗8H|�9��9$G��[m�ˑ �`c�VbY�8!��Ĳ�F��h+@���F�)����QJ�&b��&`��*D��.��!�P�� �og��F������?2���7��r��2:��m��j�>�M������aD�X��F�e6�Pe�)���~>t��u���꺺b��sHM¬�<�e�It�p�z��Kl0 >d�Pl*����"p��sG�^�L�� �����v��ˇ*]�<�4�E6h`(�y.Z�}A�5iQ�n��|�ҵ!�ԩ�<8$����,ɤ	S�p��Ll�����P�"
_��$�8�	K�1�}X�@�|_��M�B���I�7j����i� �`����� +����{H>X&�������ݟ�	�r�`8�C*�ib9-N�^z�MW�+�� �3���#0�	,����åT�Q�NL��U7d�~��F��Py��1l����HI��y	���~�PK   �x�V*�ŀ�+  �3            ��    cirkitFile.jsonPK   �x�Vs�7+5J  dK  /           ��,,  images/6c71542d-16cb-4630-930f-71c4de5e1144.pngPK   �x�V��4�� ̻ /           ���v  images/7a4be1c8-201b-41f2-b584-263fc50cb409.pngPK   �x�V]�!��	 &	 /           ���2 images/98931e0d-18f3-449f-8fca-8d5f6b2df0a7.pngPK   �x�V6�0{ { /           ��F images/c51b28eb-c857-4ce7-b81a-d633a3d7e747.pngPK   �x�V��K� 	� /           ���� images/cd1eebff-8d4c-4172-8358-6f93b12ef793.pngPK   �x�V��!�D�  Ԟ  /           ��%\ images/cf2dd1a8-295d-437f-92b8-7fcc138ae9be.pngPK   �x�VLp               ���� jsons/user_defined.jsonPK      �  ��   